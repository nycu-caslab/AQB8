
//------> /cad/mentor/Catapult/2024.1/Mgc_home/pkgs/siflibs/ccs_in_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_wait_v1 (idat, rdy, ivld, dat, irdy, vld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             rdy;
  output             ivld;
  input  [width-1:0] dat;
  input              irdy;
  input              vld;

  wire   [width-1:0] idat;
  wire               rdy;
  wire               ivld;

  localparam stallOff = 0; 
  wire                  stall_ctrl;
  assign stall_ctrl = stallOff;

  assign idat = dat;
  assign rdy = irdy && !stall_ctrl;
  assign ivld = vld && !stall_ctrl;

endmodule


//------> /cad/mentor/Catapult/2024.1/Mgc_home/pkgs/siflibs/ccs_out_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_out_wait_v1 (dat, irdy, vld, idat, rdy, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             irdy;
  output             vld;
  input  [width-1:0] idat;
  input              rdy;
  input              ivld;

  wire   [width-1:0] dat;
  wire               irdy;
  wire               vld;

  localparam stallOff = 0; 
  wire stall_ctrl;
  assign stall_ctrl = stallOff;

  assign dat = idat;
  assign irdy = rdy && !stall_ctrl;
  assign vld = ivld && !stall_ctrl;

endmodule



//------> /cad/mentor/Catapult/2024.1/Mgc_home/pkgs/siflibs/dware/ccs_dw_lp_piped_fp_recip_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - dware wrappers
//
// Copyright (c) 2021 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

// DW_lp_piped_fp_recip

//module ccs_dw_lp_piped_fp_recip_v1 (clk,rst_n,a,rnd,z,status,launch,pipe_full,pipe_ovf,accept_n,arrive,push_out_n,pipe_census);
module ccs_dw_lp_piped_fp_recip_v1 (clk,a_rst,s_rst,a,rnd,z,status,launch,pipe_full,pipe_ovf,accept_n,arrive,push_out_n,pipe_census);

  // parameters configured from C++ or hardcoded as localparam
  parameter  integer sig_width       = 23; // range 2 to 253
  parameter  integer exp_width       = 8;  // range 3 to 31
  parameter  integer ieee_compliance = 1;  // range 0 to 1
  localparam integer faithful_round  = 0;  // hardcode to 0
  localparam integer op_iso_mode     = 0;  // default
  localparam integer id_width        = 1;  // IDs not used
  parameter  integer in_reg          = 1;
  parameter  integer stages          = 4;
  parameter  integer out_reg         = 0;
  parameter  integer no_pm           = 0;
  parameter  has_rst_a               = 1;  // 1 if Catapult design uses ASync reset, 0 if Sync reset
  parameter  has_rst_s               = 0;  // Obsolete
  parameter  ph_arst                 = 0;  // Polarity of ASync reset if used
  parameter  ph_srst                 = 0;  // Polarity of Sync reset if used
  localparam rst_mode                = $unsigned(has_rst_a == 0) ? 1 : 0; // Acc to Synopsys data sheet, rst_mode=0:Async Rst; rst_mode=1:Sync Rst

  input                            clk;
  input                            a_rst;  // Async reset (has priority over sync reset)
  input                            s_rst;  // Sync reset
  input  [(sig_width+exp_width):0] a;
  input  [2:0]                     rnd;
  output [(sig_width+exp_width):0] z;
  output [7:0]                     status;
  input                            launch;
  wire   [id_width-1:0]            launch_id;
  output                           pipe_full;
  output                           pipe_ovf;
  input                            accept_n;
  output                           arrive;
  wire   [id_width-1:0]            arrive_id;
  output                           push_out_n;
  output [(((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>256)?((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>4096)?((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>16384)?((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>32768)?16:15):((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>8192)?14:13)):((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>1024)?((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>2048)?12:11):((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>512)?10:9))):((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>16)?((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>64)?((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>128)?8:7):((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>32)?6:5)):((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>4)?((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>8)?4:3):((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>2)?2:1)))))-1:0] pipe_census;
  wire                             rst_n;  // Local reset signal with polarity adjusted to be active low

  generate
  if ((has_rst_a==1)&&(ph_arst==0))
  begin: ASYNC_RESET_LOW
    assign rst_n = a_rst;
    DW_lp_piped_fp_recip #(sig_width, exp_width, ieee_compliance, 
                           faithful_round, op_iso_mode, id_width, 
                           in_reg, stages, out_reg, no_pm, rst_mode)
    U1 (.clk(clk), .rst_n(rst_n), .a(a), .rnd(rnd), .z(z), .status(status), 
          .launch(launch), .launch_id(launch_id), .pipe_full(pipe_full), .pipe_ovf(pipe_ovf),
          .accept_n(accept_n), .arrive(arrive), .arrive_id(arrive_id), .push_out_n(push_out_n), .pipe_census(pipe_census));
  end
  else if ((has_rst_a==1)&&(ph_arst==1))
  begin: ASYNC_RESET_HIGH
    assign rst_n = ~a_rst;
    DW_lp_piped_fp_recip #(sig_width, exp_width, ieee_compliance, 
                           faithful_round, op_iso_mode, id_width, 
                           in_reg, stages, out_reg, no_pm, rst_mode)
    U1 (.clk(clk), .rst_n(rst_n), .a(a), .rnd(rnd), .z(z), .status(status), 
          .launch(launch), .launch_id(launch_id), .pipe_full(pipe_full), .pipe_ovf(pipe_ovf),
          .accept_n(accept_n), .arrive(arrive), .arrive_id(arrive_id), .push_out_n(push_out_n), .pipe_census(pipe_census));
  end
  else if ((has_rst_a==0)&&(ph_srst==0))
  begin: SYNC_RESET_LOW
    assign rst_n = s_rst;
    DW_lp_piped_fp_recip #(sig_width, exp_width, ieee_compliance, 
                           faithful_round, op_iso_mode, id_width, 
                           in_reg, stages, out_reg, no_pm, rst_mode)
    U1 (.clk(clk), .rst_n(rst_n), .a(a), .rnd(rnd), .z(z), .status(status), 
          .launch(launch), .launch_id(launch_id), .pipe_full(pipe_full), .pipe_ovf(pipe_ovf),
          .accept_n(accept_n), .arrive(arrive), .arrive_id(arrive_id), .push_out_n(push_out_n), .pipe_census(pipe_census));
  end
  else if ((has_rst_a==0)&&(ph_srst==1))
  begin: SYNC_RESET_HIGH
    assign rst_n = ~s_rst;
    DW_lp_piped_fp_recip #(sig_width, exp_width, ieee_compliance, 
                           faithful_round, op_iso_mode, id_width, 
                           in_reg, stages, out_reg, no_pm, rst_mode)
    U1 (.clk(clk), .rst_n(rst_n), .a(a), .rnd(rnd), .z(z), .status(status), 
          .launch(launch), .launch_id(launch_id), .pipe_full(pipe_full), .pipe_ovf(pipe_ovf),
          .accept_n(accept_n), .arrive(arrive), .arrive_id(arrive_id), .push_out_n(push_out_n), .pipe_census(pipe_census));
  end
  endgenerate
endmodule


//------> /cad/mentor/Catapult/2024.1/Mgc_home/pkgs/siflibs/dware/ccs_dw_lp_piped_fp_add_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - dware wrappers
//
// Copyright (c) 2021 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

// DW_lp_piped_fp_add

module ccs_dw_lp_piped_fp_add_v1 (clk,a_rst,s_rst,a,b,rnd,z,status,launch,pipe_full,pipe_ovf,accept_n,arrive,push_out_n,pipe_census);
  parameter  integer sig_width       = 23; // range 2 to 253
  parameter  integer exp_width       = 8;  // range 3 to 31
  parameter  integer ieee_compliance = 1;  // range 0 to 1
  localparam integer op_iso_mode     = 0;  // hardcoded to 0
  localparam integer id_width        = 1;  // IDs not used
  parameter  integer in_reg          = 1;
  parameter  integer stages          = 4;
  parameter  integer out_reg         = 0;
  parameter  integer no_pm           = 0;
  parameter  has_rst_a               = 1;  // 1 if Catapult design uses ASync reset, 0 if Sync reset
  parameter  has_rst_s               = 0;  // Obsolete
  parameter  ph_arst                 = 0;  // Polarity of ASync reset if used
  parameter  ph_srst                 = 0;  // Polarity of Sync reset if used
  localparam rst_mode                = $unsigned(has_rst_a == 0) ? 1 : 0; // Acc to Synopsys data sheet, rst_mode=0:Async Rst; rst_mode=1:Sync Rst

  input                            clk;
  input                            a_rst;  // Async reset (has priority over sync reset)
  input                            s_rst;  // Sync reset
  input  [(sig_width+exp_width):0] a;
  input  [(sig_width+exp_width):0] b;
  input  [2:0]                     rnd;
  output [(sig_width+exp_width):0] z;
  output [7:0]                     status;
  input                            launch;
  wire   [id_width-1:0]            launch_id;
  output                           pipe_full;
  output                           pipe_ovf;
  input                            accept_n;
  output                           arrive;
  wire   [id_width-1:0]            arrive_id;
  output                           push_out_n;
  output [(((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>256)?((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>4096)?((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>16384)?((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>32768)?16:15):((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>8192)?14:13)):((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>1024)?((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>2048)?12:11):((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>512)?10:9))):((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>16)?((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>64)?((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>128)?8:7):((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>32)?6:5)):((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>4)?((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>8)?4:3):((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>2)?2:1)))))-1:0] pipe_census;
  wire                             rst_n;  // Local reset signal with polarity adjusted to be active low

  generate
  if ((has_rst_a==1)&&(ph_arst==0))
  begin: ASYNC_RESET_LOW
    assign rst_n = a_rst;
    DW_lp_piped_fp_add #(sig_width, exp_width, ieee_compliance,
        op_iso_mode, id_width,
        in_reg, stages, out_reg, no_pm, rst_mode)
      U1 (.clk(clk), .rst_n(rst_n), .a(a), .b(b), .rnd(rnd), .z(z), .status(status),
        .launch(launch), .launch_id(launch_id), .pipe_full(pipe_full), .pipe_ovf(pipe_ovf),
        .accept_n(accept_n), .arrive(arrive), .arrive_id(arrive_id), .push_out_n(push_out_n), .pipe_census(pipe_census));
  end
  else if ((has_rst_a==1)&&(ph_arst==1))
  begin: ASYNC_RESET_HIGH
    assign rst_n = ~a_rst;
    DW_lp_piped_fp_add #(sig_width, exp_width, ieee_compliance,
        op_iso_mode, id_width,
        in_reg, stages, out_reg, no_pm, rst_mode)
      U1 (.clk(clk), .rst_n(rst_n), .a(a), .b(b), .rnd(rnd), .z(z), .status(status),
        .launch(launch), .launch_id(launch_id), .pipe_full(pipe_full), .pipe_ovf(pipe_ovf),
        .accept_n(accept_n), .arrive(arrive), .arrive_id(arrive_id), .push_out_n(push_out_n), .pipe_census(pipe_census));
  end
  else if ((has_rst_a==0)&&(ph_srst==0))
  begin: SYNC_RESET_LOW
    assign rst_n = s_rst;
    DW_lp_piped_fp_add #(sig_width, exp_width, ieee_compliance,
        op_iso_mode, id_width,
        in_reg, stages, out_reg, no_pm, rst_mode)
      U1 (.clk(clk), .rst_n(rst_n), .a(a), .b(b), .rnd(rnd), .z(z), .status(status),
        .launch(launch), .launch_id(launch_id), .pipe_full(pipe_full), .pipe_ovf(pipe_ovf),
        .accept_n(accept_n), .arrive(arrive), .arrive_id(arrive_id), .push_out_n(push_out_n), .pipe_census(pipe_census));
  end
  else if ((has_rst_a==0)&&(ph_srst==1))
  begin: SYNC_RESET_HIGH
    assign rst_n = ~s_rst;
    DW_lp_piped_fp_add #(sig_width, exp_width, ieee_compliance,
        op_iso_mode, id_width,
        in_reg, stages, out_reg, no_pm, rst_mode)
      U1 (.clk(clk), .rst_n(rst_n), .a(a), .b(b), .rnd(rnd), .z(z), .status(status),
        .launch(launch), .launch_id(launch_id), .pipe_full(pipe_full), .pipe_ovf(pipe_ovf),
        .accept_n(accept_n), .arrive(arrive), .arrive_id(arrive_id), .push_out_n(push_out_n), .pipe_census(pipe_census));
  end
  endgenerate
endmodule


//------> /cad/mentor/Catapult/2024.1/Mgc_home/pkgs/siflibs/dware/ccs_dw_lp_piped_fp_mult_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - dware wrappers
//
// Copyright (c) 2021 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

// DW_lp_piped_fp_mult

module ccs_dw_lp_piped_fp_mult_v1 (clk,a_rst,s_rst,a,b,rnd,z,status,launch,pipe_full,pipe_ovf,accept_n,arrive,push_out_n,pipe_census);

  // parameters configured from C++ or hardcoded as localparam
  parameter  integer sig_width       = 23; // range 2 to 253
  parameter  integer exp_width       = 8;  // range 3 to 31
  parameter  integer ieee_compliance = 1;  // range 0 to 1
  localparam integer op_iso_mode     = 0;  // hardcode to 0
  localparam integer id_width        = 1;  // IDs not used
  parameter  integer in_reg          = 1;
  parameter  integer stages          = 4;
  parameter  integer out_reg         = 0;
  parameter  integer no_pm           = 0;
  parameter  has_rst_a               = 1;  // 1 if Catapult design uses ASync reset, 0 if Sync reset
  parameter  has_rst_s               = 0;  // Obsolete
  parameter  ph_arst                 = 0;  // Polarity of ASync reset if used
  parameter  ph_srst                 = 0;  // Polarity of Sync reset if used
  localparam rst_mode                = $unsigned(has_rst_a == 0) ? 1 : 0; // Acc to Synopsys data sheet, rst_mode=0:Async Rst; rst_mode=1:Sync Rst

  input                            clk;
  input                            a_rst;  // Async reset (has priority over sync reset)
  input                            s_rst;  // Sync reset
  input  [(sig_width+exp_width):0] a;
  input  [(sig_width+exp_width):0] b;
  input  [2:0]                     rnd;
  output [(sig_width+exp_width):0] z;
  output [7:0]                     status;
  input                            launch;
  wire   [id_width-1:0]            launch_id;
  output                           pipe_full;
  output                           pipe_ovf;
  input                            accept_n;
  output                           arrive;
  wire   [id_width-1:0]            arrive_id;
  output                           push_out_n;
  output [(((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>256)?((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>4096)?((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>16384)?((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>32768)?16:15):((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>8192)?14:13)):((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>1024)?((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>2048)?12:11):((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>512)?10:9))):((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>16)?((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>64)?((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>128)?8:7):((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>32)?6:5)):((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>4)?((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>8)?4:3):((((((in_reg+(stages-1)+out_reg) >= 1) ? (in_reg+(stages-1)+out_reg) : 1)+1)>2)?2:1)))))-1:0] pipe_census;
  wire                             rst_n;  // Local reset signal with polarity adjusted to be active low

  generate
  if ((has_rst_a==1)&&(ph_arst==0))
  begin: ASYNC_RESET_LOW
    assign rst_n = a_rst;
    DW_lp_piped_fp_mult #(sig_width, exp_width, ieee_compliance,
        op_iso_mode, id_width,
        in_reg, stages, out_reg, no_pm, rst_mode)
      U1 (.clk(clk), .rst_n(rst_n), .a(a), .b(b), .rnd(rnd), .z(z), .status(status),
        .launch(launch), .launch_id(launch_id), .pipe_full(pipe_full), .pipe_ovf(pipe_ovf),
        .accept_n(accept_n), .arrive(arrive), .arrive_id(arrive_id), .push_out_n(push_out_n), .pipe_census(pipe_census));
  end
  else if ((has_rst_a==1)&&(ph_arst==1))
  begin: ASYNC_RESET_HIGH
    assign rst_n = ~a_rst;
    DW_lp_piped_fp_mult #(sig_width, exp_width, ieee_compliance,
        op_iso_mode, id_width,
        in_reg, stages, out_reg, no_pm, rst_mode)
      U1 (.clk(clk), .rst_n(rst_n), .a(a), .b(b), .rnd(rnd), .z(z), .status(status),
        .launch(launch), .launch_id(launch_id), .pipe_full(pipe_full), .pipe_ovf(pipe_ovf),
        .accept_n(accept_n), .arrive(arrive), .arrive_id(arrive_id), .push_out_n(push_out_n), .pipe_census(pipe_census));
  end
  else if ((has_rst_a==0)&&(ph_srst==0))
  begin: SYNC_RESET_LOW
    assign rst_n = s_rst;
    DW_lp_piped_fp_mult #(sig_width, exp_width, ieee_compliance,
        op_iso_mode, id_width,
        in_reg, stages, out_reg, no_pm, rst_mode)
      U1 (.clk(clk), .rst_n(rst_n), .a(a), .b(b), .rnd(rnd), .z(z), .status(status),
        .launch(launch), .launch_id(launch_id), .pipe_full(pipe_full), .pipe_ovf(pipe_ovf),
        .accept_n(accept_n), .arrive(arrive), .arrive_id(arrive_id), .push_out_n(push_out_n), .pipe_census(pipe_census));
  end
  else if ((has_rst_a==0)&&(ph_srst==1))
  begin: SYNC_RESET_HIGH
    assign rst_n = ~s_rst;
    DW_lp_piped_fp_mult #(sig_width, exp_width, ieee_compliance,
        op_iso_mode, id_width,
        in_reg, stages, out_reg, no_pm, rst_mode)
      U1 (.clk(clk), .rst_n(rst_n), .a(a), .b(b), .rnd(rnd), .z(z), .status(status),
        .launch(launch), .launch_id(launch_id), .pipe_full(pipe_full), .pipe_ovf(pipe_ovf),
        .accept_n(accept_n), .arrive(arrive), .arrive_id(arrive_id), .push_out_n(push_out_n), .pipe_census(pipe_census));
  end
  endgenerate
endmodule


//------> /cad/mentor/Catapult/2024.1/Mgc_home/pkgs/siflibs/dware/ccs_dw_fp_cmp_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - dware wrappers
//
// Copyright (c) 2021 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

// DW_fp_cmp

module ccs_dw_fp_cmp_v1 (a, b, zctr, aeqb, altb, agtb, unordered, z0, z1, status0, status1);
  parameter  integer sig_width = 23;      // range 2 to 253
  parameter  integer exp_width = 8;       // range 3 to 31
  parameter  integer ieee_compliance = 0; // range 0 to 1
  input  [sig_width + exp_width:0] a;
  input  [sig_width + exp_width:0] b;
  input  zctr;
  output aeqb, altb, agtb, unordered;
  output [sig_width + exp_width:0] z0, z1;
  output [7:0] status0, status1;

  DW_fp_cmp #(sig_width,exp_width,ieee_compliance)
    U1 (.a(a), .b(b), .zctr(zctr), .aeqb(aeqb), .altb(altb), .agtb(agtb), .unordered(unordered), .z0(z0), .z1(z1), .status0(status0), .status1(status1));
endmodule

//------> /cad/mentor/Catapult/2024.1/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.v 
module mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ../td_ccore_solutions/leading_sign_8_0_1_0_8d285dc35b24d6e9e4ec5943bd36901f5975_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   lashhw@localhost.localdomain
//  Generated date: Fri Jan 31 20:29:12 2025
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    leading_sign_8_0_1_0
// ------------------------------------------------------------------


module leading_sign_8_0_1_0 (
  mantissa, rtn
);
  input [7:0] mantissa;
  output [3:0] rtn;


  // Interconnect Declarations
  wire ac_private_LeadingSignConstrained_true_false_val_133_8_false_all_sign_wrs_c_6_2_sdt_2;
  wire ac_private_LeadingSignConstrained_true_false_val_133_8_false_all_sign_wrs_c_20_3_sdt_3;
  wire ac_private_LeadingSignConstrained_true_false_val_133_8_false_all_sign_wrs_c_6_2_sdt_1;
  wire ac_private_LeadingSignConstrained_true_false_val_133_8_false_all_sign_wrs_c_14_2_sdt_1;
  wire c_h_1_2;

  wire[2:0] ac_private_LeadingSignConstrained_true_false_val_133_8_false_all_sign_ac_private_LeadingSignConstrained_true_false_val_133_8_false_all_sign_and_nl;
  wire ac_private_LeadingSignConstrained_true_false_val_133_8_false_all_sign_and_23_nl;
  wire ac_private_LeadingSignConstrained_true_false_val_133_8_false_all_sign_and_21_nl;
  wire ac_private_LeadingSignConstrained_true_false_val_133_8_false_all_sign_not_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ac_private_LeadingSignConstrained_true_false_val_133_8_false_all_sign_wrs_c_6_2_sdt_2
      = ~((mantissa[5:4]!=2'b00));
  assign ac_private_LeadingSignConstrained_true_false_val_133_8_false_all_sign_wrs_c_6_2_sdt_1
      = ~((mantissa[7:6]!=2'b00));
  assign ac_private_LeadingSignConstrained_true_false_val_133_8_false_all_sign_wrs_c_14_2_sdt_1
      = ~((mantissa[3:2]!=2'b00));
  assign c_h_1_2 = ac_private_LeadingSignConstrained_true_false_val_133_8_false_all_sign_wrs_c_6_2_sdt_1
      & ac_private_LeadingSignConstrained_true_false_val_133_8_false_all_sign_wrs_c_6_2_sdt_2;
  assign ac_private_LeadingSignConstrained_true_false_val_133_8_false_all_sign_wrs_c_20_3_sdt_3
      = (mantissa[1:0]==2'b00) & ac_private_LeadingSignConstrained_true_false_val_133_8_false_all_sign_wrs_c_14_2_sdt_1
      & c_h_1_2;
  assign ac_private_LeadingSignConstrained_true_false_val_133_8_false_all_sign_and_23_nl
      = ac_private_LeadingSignConstrained_true_false_val_133_8_false_all_sign_wrs_c_6_2_sdt_1
      & (ac_private_LeadingSignConstrained_true_false_val_133_8_false_all_sign_wrs_c_14_2_sdt_1
      | (~ ac_private_LeadingSignConstrained_true_false_val_133_8_false_all_sign_wrs_c_6_2_sdt_2));
  assign ac_private_LeadingSignConstrained_true_false_val_133_8_false_all_sign_and_21_nl
      = (~((mantissa[7]) | (~((mantissa[6:5]!=2'b01))))) & (~(((mantissa[3]) | (~((mantissa[2:1]!=2'b01))))
      & c_h_1_2));
  assign ac_private_LeadingSignConstrained_true_false_val_133_8_false_all_sign_not_nl
      = ~ ac_private_LeadingSignConstrained_true_false_val_133_8_false_all_sign_wrs_c_20_3_sdt_3;
  assign ac_private_LeadingSignConstrained_true_false_val_133_8_false_all_sign_ac_private_LeadingSignConstrained_true_false_val_133_8_false_all_sign_and_nl
      = MUX_v_3_2_2(3'b000, ({c_h_1_2 , ac_private_LeadingSignConstrained_true_false_val_133_8_false_all_sign_and_23_nl
      , ac_private_LeadingSignConstrained_true_false_val_133_8_false_all_sign_and_21_nl}),
      ac_private_LeadingSignConstrained_true_false_val_133_8_false_all_sign_not_nl);
  assign rtn = {ac_private_LeadingSignConstrained_true_false_val_133_8_false_all_sign_wrs_c_20_3_sdt_3
      , ac_private_LeadingSignConstrained_true_false_val_133_8_false_all_sign_ac_private_LeadingSignConstrained_true_false_val_133_8_false_all_sign_and_nl};

  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input  sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction

endmodule




//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2024.1/1091966 Production Release
//  HLS Date:       Wed Feb 14 09:07:18 PST 2024
// 
//  Generated by:   lashhw@localhost.localdomain
//  Generated date: Fri Jan 31 22:39:30 2025
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    init_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module init_core_core_fsm (
  clk, arst_n, core_wen, fsm_output
);
  input clk;
  input arst_n;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for init_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg  state_var;
  reg  state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : init_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_staller
// ------------------------------------------------------------------


module init_core_staller (
  clk, arst_n, core_wen, core_wten, init_req_stream_rsci_wen_comp, trv_req_stream_rsci_wen_comp,
      core_flen_unreg
);
  input clk;
  input arst_n;
  output core_wen;
  output core_wten;
  input init_req_stream_rsci_wen_comp;
  input trv_req_stream_rsci_wen_comp;
  input core_flen_unreg;


  // Interconnect Declarations
  reg core_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign core_wen = init_req_stream_rsci_wen_comp & trv_req_stream_rsci_wen_comp
      & (~ core_flen_unreg);
  assign core_wten = core_wten_reg;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      core_wten_reg <= 1'b0;
    end
    else begin
      core_wten_reg <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_2_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_dp_2
// ------------------------------------------------------------------


module init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_2_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_dp_2
    (
  clk, arst_n, ccs_lp_piped_fp_recip_23_8_0_cmp_2_bawt, ccs_lp_piped_fp_recip_23_8_0_cmp_2_z_mxwt,
      ccs_lp_piped_fp_recip_23_8_0_cmp_2_biwt, ccs_lp_piped_fp_recip_23_8_0_cmp_2_bdwt,
      ccs_lp_piped_fp_recip_23_8_0_cmp_2_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_recip_23_8_0_cmp_2_bawt;
  output [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_2_z_mxwt;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_2_biwt;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_2_bdwt;
  input [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_2_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_recip_23_8_0_cmp_2_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_recip_23_8_0_cmp_2_bcwt;
  reg [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_2_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_2_z_bfwt_1;

  wire[1:0] lp_piped_fp_recip_AC_RND_CONV_0_32_8_1_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_recip_AC_RND_CONV_0_32_8_1_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_recip_23_8_0_cmp_2_bawt = ccs_lp_piped_fp_recip_23_8_0_cmp_2_biwt
      | (ccs_lp_piped_fp_recip_23_8_0_cmp_2_bcwt!=2'b00);
  assign ccs_lp_piped_fp_recip_23_8_0_cmp_2_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_recip_23_8_0_cmp_2_z,
      ccs_lp_piped_fp_recip_23_8_0_cmp_2_z_bfwt, ccs_lp_piped_fp_recip_23_8_0_cmp_2_z_bfwt_1,
      ccs_lp_piped_fp_recip_23_8_0_cmp_2_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_recip_23_8_0_cmp_2_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_recip_23_8_0_cmp_2_bcwt <= nl_ccs_lp_piped_fp_recip_23_8_0_cmp_2_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_recip_23_8_0_cmp_2_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_recip_23_8_0_cmp_2_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_recip_23_8_0_cmp_2_biwt ) begin
      ccs_lp_piped_fp_recip_23_8_0_cmp_2_z_bfwt <= ccs_lp_piped_fp_recip_23_8_0_cmp_2_z;
      ccs_lp_piped_fp_recip_23_8_0_cmp_2_z_bfwt_1 <= ccs_lp_piped_fp_recip_23_8_0_cmp_2_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_recip_AC_RND_CONV_0_32_8_1_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_recip_23_8_0_cmp_2_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_recip_23_8_0_cmp_2_biwt);
  assign lp_piped_fp_recip_AC_RND_CONV_0_32_8_1_acc_1_nl = nl_lp_piped_fp_recip_AC_RND_CONV_0_32_8_1_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_recip_23_8_0_cmp_2_bcwt  = lp_piped_fp_recip_AC_RND_CONV_0_32_8_1_acc_1_nl
      + ccs_lp_piped_fp_recip_23_8_0_cmp_2_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_2_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_ctrl_2
// ------------------------------------------------------------------


module init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_2_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_ctrl_2
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_recip_23_8_0_cmp_2_oswt_unreg,
      ccs_lp_piped_fp_recip_23_8_0_cmp_2_iswt1, ccs_lp_piped_fp_recip_23_8_0_cmp_2_biwt,
      ccs_lp_piped_fp_recip_23_8_0_cmp_2_bdwt, ccs_lp_piped_fp_recip_23_8_0_cmp_2_launch_core_sct,
      ccs_lp_piped_fp_recip_23_8_0_cmp_2_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_2_oswt_unreg;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_2_iswt1;
  output ccs_lp_piped_fp_recip_23_8_0_cmp_2_biwt;
  output ccs_lp_piped_fp_recip_23_8_0_cmp_2_bdwt;
  output ccs_lp_piped_fp_recip_23_8_0_cmp_2_launch_core_sct;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_2_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_recip_23_8_0_cmp_2_cs_lp_piped_fp_recip_23_8_0_cmp_2_pdswt0;
  reg [1:0] ccs_lp_piped_fp_recip_23_8_0_cmp_2_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_recip_23_8_0_cmp_2_icwt;

  wire[1:0] lp_piped_fp_recip_AC_RND_CONV_0_32_8_1_acc_nl;
  wire[2:0] nl_lp_piped_fp_recip_AC_RND_CONV_0_32_8_1_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_recip_23_8_0_cmp_2_bdwt = ccs_lp_piped_fp_recip_23_8_0_cmp_2_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_recip_23_8_0_cmp_2_biwt = ccs_lp_piped_fp_recip_23_8_0_cmp_2_cs_lp_piped_fp_recip_23_8_0_cmp_2_pdswt0
      | (ccs_lp_piped_fp_recip_23_8_0_cmp_2_icwt!=2'b00);
  assign ccs_lp_piped_fp_recip_23_8_0_cmp_2_launch_core_sct = core_wen & ccs_lp_piped_fp_recip_23_8_0_cmp_2_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_recip_23_8_0_cmp_2_cs_lp_piped_fp_recip_23_8_0_cmp_2_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_recip_23_8_0_cmp_2_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_recip_23_8_0_cmp_2_cs_lp_piped_fp_recip_23_8_0_cmp_2_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_recip_23_8_0_cmp_2_iswt1;
      ccs_lp_piped_fp_recip_23_8_0_cmp_2_icwt <= nl_ccs_lp_piped_fp_recip_23_8_0_cmp_2_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_recip_AC_RND_CONV_0_32_8_1_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_recip_23_8_0_cmp_2_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_recip_23_8_0_cmp_2_cs_lp_piped_fp_recip_23_8_0_cmp_2_pdswt0);
  assign lp_piped_fp_recip_AC_RND_CONV_0_32_8_1_acc_nl = nl_lp_piped_fp_recip_AC_RND_CONV_0_32_8_1_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_recip_23_8_0_cmp_2_icwt  = lp_piped_fp_recip_AC_RND_CONV_0_32_8_1_acc_nl
      + ccs_lp_piped_fp_recip_23_8_0_cmp_2_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_1_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_dp_1
// ------------------------------------------------------------------


module init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_1_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_dp_1
    (
  clk, arst_n, ccs_lp_piped_fp_recip_23_8_0_cmp_1_bawt, ccs_lp_piped_fp_recip_23_8_0_cmp_1_z_mxwt,
      ccs_lp_piped_fp_recip_23_8_0_cmp_1_biwt, ccs_lp_piped_fp_recip_23_8_0_cmp_1_bdwt,
      ccs_lp_piped_fp_recip_23_8_0_cmp_1_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_recip_23_8_0_cmp_1_bawt;
  output [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_1_z_mxwt;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_1_biwt;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_1_bdwt;
  input [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_1_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_recip_23_8_0_cmp_1_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_recip_23_8_0_cmp_1_bcwt;
  reg [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_1_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_1_z_bfwt_1;

  wire[1:0] lp_piped_fp_recip_AC_RND_CONV_0_32_8_2_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_recip_AC_RND_CONV_0_32_8_2_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_recip_23_8_0_cmp_1_bawt = ccs_lp_piped_fp_recip_23_8_0_cmp_1_biwt
      | (ccs_lp_piped_fp_recip_23_8_0_cmp_1_bcwt!=2'b00);
  assign ccs_lp_piped_fp_recip_23_8_0_cmp_1_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_recip_23_8_0_cmp_1_z,
      ccs_lp_piped_fp_recip_23_8_0_cmp_1_z_bfwt, ccs_lp_piped_fp_recip_23_8_0_cmp_1_z_bfwt_1,
      ccs_lp_piped_fp_recip_23_8_0_cmp_1_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_recip_23_8_0_cmp_1_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_recip_23_8_0_cmp_1_bcwt <= nl_ccs_lp_piped_fp_recip_23_8_0_cmp_1_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_recip_23_8_0_cmp_1_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_recip_23_8_0_cmp_1_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_recip_23_8_0_cmp_1_biwt ) begin
      ccs_lp_piped_fp_recip_23_8_0_cmp_1_z_bfwt <= ccs_lp_piped_fp_recip_23_8_0_cmp_1_z;
      ccs_lp_piped_fp_recip_23_8_0_cmp_1_z_bfwt_1 <= ccs_lp_piped_fp_recip_23_8_0_cmp_1_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_recip_AC_RND_CONV_0_32_8_2_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_recip_23_8_0_cmp_1_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_recip_23_8_0_cmp_1_biwt);
  assign lp_piped_fp_recip_AC_RND_CONV_0_32_8_2_acc_1_nl = nl_lp_piped_fp_recip_AC_RND_CONV_0_32_8_2_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_recip_23_8_0_cmp_1_bcwt  = lp_piped_fp_recip_AC_RND_CONV_0_32_8_2_acc_1_nl
      + ccs_lp_piped_fp_recip_23_8_0_cmp_1_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_1_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_ctrl_1
// ------------------------------------------------------------------


module init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_1_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_ctrl_1
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_recip_23_8_0_cmp_1_oswt_unreg,
      ccs_lp_piped_fp_recip_23_8_0_cmp_1_iswt1, ccs_lp_piped_fp_recip_23_8_0_cmp_1_biwt,
      ccs_lp_piped_fp_recip_23_8_0_cmp_1_bdwt, ccs_lp_piped_fp_recip_23_8_0_cmp_1_launch_core_sct,
      ccs_lp_piped_fp_recip_23_8_0_cmp_1_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_1_oswt_unreg;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_1_iswt1;
  output ccs_lp_piped_fp_recip_23_8_0_cmp_1_biwt;
  output ccs_lp_piped_fp_recip_23_8_0_cmp_1_bdwt;
  output ccs_lp_piped_fp_recip_23_8_0_cmp_1_launch_core_sct;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_1_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_recip_23_8_0_cmp_1_cs_lp_piped_fp_recip_23_8_0_cmp_1_pdswt0;
  reg [1:0] ccs_lp_piped_fp_recip_23_8_0_cmp_1_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_recip_23_8_0_cmp_1_icwt;

  wire[1:0] lp_piped_fp_recip_AC_RND_CONV_0_32_8_2_acc_nl;
  wire[2:0] nl_lp_piped_fp_recip_AC_RND_CONV_0_32_8_2_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_recip_23_8_0_cmp_1_bdwt = ccs_lp_piped_fp_recip_23_8_0_cmp_1_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_recip_23_8_0_cmp_1_biwt = ccs_lp_piped_fp_recip_23_8_0_cmp_1_cs_lp_piped_fp_recip_23_8_0_cmp_1_pdswt0
      | (ccs_lp_piped_fp_recip_23_8_0_cmp_1_icwt!=2'b00);
  assign ccs_lp_piped_fp_recip_23_8_0_cmp_1_launch_core_sct = core_wen & ccs_lp_piped_fp_recip_23_8_0_cmp_1_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_recip_23_8_0_cmp_1_cs_lp_piped_fp_recip_23_8_0_cmp_1_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_recip_23_8_0_cmp_1_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_recip_23_8_0_cmp_1_cs_lp_piped_fp_recip_23_8_0_cmp_1_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_recip_23_8_0_cmp_1_iswt1;
      ccs_lp_piped_fp_recip_23_8_0_cmp_1_icwt <= nl_ccs_lp_piped_fp_recip_23_8_0_cmp_1_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_recip_AC_RND_CONV_0_32_8_2_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_recip_23_8_0_cmp_1_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_recip_23_8_0_cmp_1_cs_lp_piped_fp_recip_23_8_0_cmp_1_pdswt0);
  assign lp_piped_fp_recip_AC_RND_CONV_0_32_8_2_acc_nl = nl_lp_piped_fp_recip_AC_RND_CONV_0_32_8_2_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_recip_23_8_0_cmp_1_icwt  = lp_piped_fp_recip_AC_RND_CONV_0_32_8_2_acc_nl
      + ccs_lp_piped_fp_recip_23_8_0_cmp_1_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_dp
// ------------------------------------------------------------------


module init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_dp
    (
  clk, arst_n, ccs_lp_piped_fp_recip_23_8_0_cmp_bawt, ccs_lp_piped_fp_recip_23_8_0_cmp_z_mxwt,
      ccs_lp_piped_fp_recip_23_8_0_cmp_biwt, ccs_lp_piped_fp_recip_23_8_0_cmp_bdwt,
      ccs_lp_piped_fp_recip_23_8_0_cmp_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_recip_23_8_0_cmp_bawt;
  output [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_z_mxwt;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_biwt;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_bdwt;
  input [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_recip_23_8_0_cmp_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_recip_23_8_0_cmp_bcwt;
  reg [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_z_bfwt_1;

  wire[1:0] lp_piped_fp_recip_AC_RND_CONV_0_32_8_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_recip_AC_RND_CONV_0_32_8_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_recip_23_8_0_cmp_bawt = ccs_lp_piped_fp_recip_23_8_0_cmp_biwt
      | (ccs_lp_piped_fp_recip_23_8_0_cmp_bcwt!=2'b00);
  assign ccs_lp_piped_fp_recip_23_8_0_cmp_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_recip_23_8_0_cmp_z,
      ccs_lp_piped_fp_recip_23_8_0_cmp_z_bfwt, ccs_lp_piped_fp_recip_23_8_0_cmp_z_bfwt_1,
      ccs_lp_piped_fp_recip_23_8_0_cmp_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_recip_23_8_0_cmp_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_recip_23_8_0_cmp_bcwt <= nl_ccs_lp_piped_fp_recip_23_8_0_cmp_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_recip_23_8_0_cmp_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_recip_23_8_0_cmp_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_recip_23_8_0_cmp_biwt ) begin
      ccs_lp_piped_fp_recip_23_8_0_cmp_z_bfwt <= ccs_lp_piped_fp_recip_23_8_0_cmp_z;
      ccs_lp_piped_fp_recip_23_8_0_cmp_z_bfwt_1 <= ccs_lp_piped_fp_recip_23_8_0_cmp_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_recip_AC_RND_CONV_0_32_8_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_recip_23_8_0_cmp_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_recip_23_8_0_cmp_biwt);
  assign lp_piped_fp_recip_AC_RND_CONV_0_32_8_acc_1_nl = nl_lp_piped_fp_recip_AC_RND_CONV_0_32_8_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_recip_23_8_0_cmp_bcwt  = lp_piped_fp_recip_AC_RND_CONV_0_32_8_acc_1_nl
      + ccs_lp_piped_fp_recip_23_8_0_cmp_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_ctrl
// ------------------------------------------------------------------


module init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_ctrl
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_recip_23_8_0_cmp_oswt_unreg,
      ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1, ccs_lp_piped_fp_recip_23_8_0_cmp_biwt,
      ccs_lp_piped_fp_recip_23_8_0_cmp_bdwt, ccs_lp_piped_fp_recip_23_8_0_cmp_launch_core_sct,
      ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_oswt_unreg;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1;
  output ccs_lp_piped_fp_recip_23_8_0_cmp_biwt;
  output ccs_lp_piped_fp_recip_23_8_0_cmp_bdwt;
  output ccs_lp_piped_fp_recip_23_8_0_cmp_launch_core_sct;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_recip_23_8_0_cmp_cs_lp_piped_fp_recip_23_8_0_cmp_pdswt0;
  reg [1:0] ccs_lp_piped_fp_recip_23_8_0_cmp_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_recip_23_8_0_cmp_icwt;

  wire[1:0] lp_piped_fp_recip_AC_RND_CONV_0_32_8_acc_nl;
  wire[2:0] nl_lp_piped_fp_recip_AC_RND_CONV_0_32_8_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_recip_23_8_0_cmp_bdwt = ccs_lp_piped_fp_recip_23_8_0_cmp_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_recip_23_8_0_cmp_biwt = ccs_lp_piped_fp_recip_23_8_0_cmp_cs_lp_piped_fp_recip_23_8_0_cmp_pdswt0
      | (ccs_lp_piped_fp_recip_23_8_0_cmp_icwt!=2'b00);
  assign ccs_lp_piped_fp_recip_23_8_0_cmp_launch_core_sct = core_wen & ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_recip_23_8_0_cmp_cs_lp_piped_fp_recip_23_8_0_cmp_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_recip_23_8_0_cmp_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_recip_23_8_0_cmp_cs_lp_piped_fp_recip_23_8_0_cmp_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1;
      ccs_lp_piped_fp_recip_23_8_0_cmp_icwt <= nl_ccs_lp_piped_fp_recip_23_8_0_cmp_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_recip_AC_RND_CONV_0_32_8_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_recip_23_8_0_cmp_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_recip_23_8_0_cmp_cs_lp_piped_fp_recip_23_8_0_cmp_pdswt0);
  assign lp_piped_fp_recip_AC_RND_CONV_0_32_8_acc_nl = nl_lp_piped_fp_recip_AC_RND_CONV_0_32_8_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_recip_23_8_0_cmp_icwt  = lp_piped_fp_recip_AC_RND_CONV_0_32_8_acc_nl
      + ccs_lp_piped_fp_recip_23_8_0_cmp_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_2
// ------------------------------------------------------------------


module init_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_2
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_2_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_2_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_2_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_2_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_2_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_2_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_2_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_2_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_2_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_2_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_2_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_2_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_2_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_2_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_2_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_2_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_2_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_2_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_2
// ------------------------------------------------------------------


module init_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_2
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_2_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_2_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_2_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_2_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_2_cs_lp_piped_fp_add_23_8_0_cmp_2_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_2_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_2_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_2_cs_lp_piped_fp_add_23_8_0_cmp_2_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_2_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_2_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_2_cs_lp_piped_fp_add_23_8_0_cmp_2_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_2_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_2_cs_lp_piped_fp_add_23_8_0_cmp_2_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_2_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_2_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_2_cs_lp_piped_fp_add_23_8_0_cmp_2_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_2_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_2_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_1
// ------------------------------------------------------------------


module init_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_1
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_1_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_1_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_1_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_1_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_1_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_1_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_1_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_1_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_1_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_1_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_1_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_1_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_1_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_1_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_1_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_1_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_1_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_1_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_1
// ------------------------------------------------------------------


module init_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_1
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_1_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_1_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_1_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_1_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_1_cs_lp_piped_fp_add_23_8_0_cmp_1_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_1_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_1_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_1_cs_lp_piped_fp_add_23_8_0_cmp_1_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_1_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_1_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_1_cs_lp_piped_fp_add_23_8_0_cmp_1_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_1_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_1_cs_lp_piped_fp_add_23_8_0_cmp_1_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_1_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_1_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_1_cs_lp_piped_fp_add_23_8_0_cmp_1_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_1_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_1_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_ccs_lp_piped_fp_add_23_8_0_cmp_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp
// ------------------------------------------------------------------


module init_core_ccs_lp_piped_fp_add_23_8_0_cmp_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_ccs_lp_piped_fp_add_23_8_0_cmp_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl
// ------------------------------------------------------------------


module init_core_ccs_lp_piped_fp_add_23_8_0_cmp_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_oswt_unreg, ccs_lp_piped_fp_add_23_8_0_cmp_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_cs_lp_piped_fp_add_23_8_0_cmp_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_cs_lp_piped_fp_add_23_8_0_cmp_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_cs_lp_piped_fp_add_23_8_0_cmp_pdswt0 <= 1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_cs_lp_piped_fp_add_23_8_0_cmp_pdswt0 <= (~ core_wten)
          & ccs_lp_piped_fp_add_23_8_0_cmp_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_cs_lp_piped_fp_add_23_8_0_cmp_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_2
// ------------------------------------------------------------------


module init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_2
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_2_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_2_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_2_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_2_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_2_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_2_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_2_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_2
// ------------------------------------------------------------------


module init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_2
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_2_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_2_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_2_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_2_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_2_cs_lp_piped_fp_mult_23_8_0_cmp_2_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_2_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_2_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_2_cs_lp_piped_fp_mult_23_8_0_cmp_2_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_2_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_2_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_cs_lp_piped_fp_mult_23_8_0_cmp_2_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_cs_lp_piped_fp_mult_23_8_0_cmp_2_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_2_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_2_cs_lp_piped_fp_mult_23_8_0_cmp_2_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_2_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_2_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_1
// ------------------------------------------------------------------


module init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_1
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_1_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_1_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_1_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_1_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_1_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_1_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_1_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_1
// ------------------------------------------------------------------


module init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_1
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_1_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_1_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_1_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_1_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_1_cs_lp_piped_fp_mult_23_8_0_cmp_1_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_1_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_1_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_1_cs_lp_piped_fp_mult_23_8_0_cmp_1_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_1_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_1_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_cs_lp_piped_fp_mult_23_8_0_cmp_1_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_cs_lp_piped_fp_mult_23_8_0_cmp_1_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_1_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_1_cs_lp_piped_fp_mult_23_8_0_cmp_1_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_1_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_1_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp
// ------------------------------------------------------------------


module init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl
// ------------------------------------------------------------------


module init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_oswt_unreg, ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_launch_core_sct, ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_cs_lp_piped_fp_mult_23_8_0_cmp_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_cs_lp_piped_fp_mult_23_8_0_cmp_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_cs_lp_piped_fp_mult_23_8_0_cmp_pdswt0 <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_cs_lp_piped_fp_mult_23_8_0_cmp_pdswt0 <= (~
          core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_cs_lp_piped_fp_mult_23_8_0_cmp_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_trv_req_stream_rsci_trv_req_stream_wait_dp
// ------------------------------------------------------------------


module init_core_trv_req_stream_rsci_trv_req_stream_wait_dp (
  clk, arst_n, trv_req_stream_rsci_oswt_unreg, trv_req_stream_rsci_bawt, trv_req_stream_rsci_wen_comp,
      trv_req_stream_rsci_biwt, trv_req_stream_rsci_bdwt, trv_req_stream_rsci_bcwt
);
  input clk;
  input arst_n;
  input trv_req_stream_rsci_oswt_unreg;
  output trv_req_stream_rsci_bawt;
  output trv_req_stream_rsci_wen_comp;
  input trv_req_stream_rsci_biwt;
  input trv_req_stream_rsci_bdwt;
  output trv_req_stream_rsci_bcwt;
  reg trv_req_stream_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign trv_req_stream_rsci_bawt = trv_req_stream_rsci_biwt | trv_req_stream_rsci_bcwt;
  assign trv_req_stream_rsci_wen_comp = (~ trv_req_stream_rsci_oswt_unreg) | trv_req_stream_rsci_bawt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      trv_req_stream_rsci_bcwt <= 1'b0;
    end
    else begin
      trv_req_stream_rsci_bcwt <= ~((~(trv_req_stream_rsci_bcwt | trv_req_stream_rsci_biwt))
          | trv_req_stream_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_trv_req_stream_rsci_trv_req_stream_wait_ctrl
// ------------------------------------------------------------------


module init_core_trv_req_stream_rsci_trv_req_stream_wait_ctrl (
  core_wen, trv_req_stream_rsci_oswt_unreg, trv_req_stream_rsci_iswt0, trv_req_stream_rsci_biwt,
      trv_req_stream_rsci_bdwt, trv_req_stream_rsci_bcwt, trv_req_stream_rsci_irdy,
      trv_req_stream_rsci_ivld_core_sct
);
  input core_wen;
  input trv_req_stream_rsci_oswt_unreg;
  input trv_req_stream_rsci_iswt0;
  output trv_req_stream_rsci_biwt;
  output trv_req_stream_rsci_bdwt;
  input trv_req_stream_rsci_bcwt;
  input trv_req_stream_rsci_irdy;
  output trv_req_stream_rsci_ivld_core_sct;


  // Interconnect Declarations
  wire trv_req_stream_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign trv_req_stream_rsci_bdwt = trv_req_stream_rsci_oswt_unreg & core_wen;
  assign trv_req_stream_rsci_biwt = trv_req_stream_rsci_ogwt & trv_req_stream_rsci_irdy;
  assign trv_req_stream_rsci_ogwt = trv_req_stream_rsci_iswt0 & (~ trv_req_stream_rsci_bcwt);
  assign trv_req_stream_rsci_ivld_core_sct = trv_req_stream_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_init_req_stream_rsci_init_req_stream_wait_dp
// ------------------------------------------------------------------


module init_core_init_req_stream_rsci_init_req_stream_wait_dp (
  clk, arst_n, init_req_stream_rsci_oswt_unreg, init_req_stream_rsci_bawt, init_req_stream_rsci_wen_comp,
      init_req_stream_rsci_idat_mxwt, init_req_stream_rsci_biwt, init_req_stream_rsci_bdwt,
      init_req_stream_rsci_bcwt, init_req_stream_rsci_idat
);
  input clk;
  input arst_n;
  input init_req_stream_rsci_oswt_unreg;
  output init_req_stream_rsci_bawt;
  output init_req_stream_rsci_wen_comp;
  output [361:0] init_req_stream_rsci_idat_mxwt;
  input init_req_stream_rsci_biwt;
  input init_req_stream_rsci_bdwt;
  output init_req_stream_rsci_bcwt;
  reg init_req_stream_rsci_bcwt;
  input [361:0] init_req_stream_rsci_idat;


  // Interconnect Declarations
  reg [361:0] init_req_stream_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign init_req_stream_rsci_bawt = init_req_stream_rsci_biwt | init_req_stream_rsci_bcwt;
  assign init_req_stream_rsci_wen_comp = (~ init_req_stream_rsci_oswt_unreg) | init_req_stream_rsci_bawt;
  assign init_req_stream_rsci_idat_mxwt = MUX_v_362_2_2(init_req_stream_rsci_idat,
      init_req_stream_rsci_idat_bfwt, init_req_stream_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      init_req_stream_rsci_bcwt <= 1'b0;
    end
    else begin
      init_req_stream_rsci_bcwt <= ~((~(init_req_stream_rsci_bcwt | init_req_stream_rsci_biwt))
          | init_req_stream_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      init_req_stream_rsci_idat_bfwt <= 362'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( init_req_stream_rsci_biwt ) begin
      init_req_stream_rsci_idat_bfwt <= init_req_stream_rsci_idat;
    end
  end

  function automatic [361:0] MUX_v_362_2_2;
    input [361:0] input_0;
    input [361:0] input_1;
    input  sel;
    reg [361:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_362_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_init_req_stream_rsci_init_req_stream_wait_ctrl
// ------------------------------------------------------------------


module init_core_init_req_stream_rsci_init_req_stream_wait_ctrl (
  core_wen, init_req_stream_rsci_oswt_unreg, init_req_stream_rsci_iswt0, init_req_stream_rsci_biwt,
      init_req_stream_rsci_bdwt, init_req_stream_rsci_bcwt, init_req_stream_rsci_irdy_core_sct,
      init_req_stream_rsci_ivld
);
  input core_wen;
  input init_req_stream_rsci_oswt_unreg;
  input init_req_stream_rsci_iswt0;
  output init_req_stream_rsci_biwt;
  output init_req_stream_rsci_bdwt;
  input init_req_stream_rsci_bcwt;
  output init_req_stream_rsci_irdy_core_sct;
  input init_req_stream_rsci_ivld;


  // Interconnect Declarations
  wire init_req_stream_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign init_req_stream_rsci_bdwt = init_req_stream_rsci_oswt_unreg & core_wen;
  assign init_req_stream_rsci_biwt = init_req_stream_rsci_ogwt & init_req_stream_rsci_ivld;
  assign init_req_stream_rsci_ogwt = init_req_stream_rsci_iswt0 & (~ init_req_stream_rsci_bcwt);
  assign init_req_stream_rsci_irdy_core_sct = init_req_stream_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module bbox_core_core_fsm (
  clk, arst_n, core_wen, fsm_output
);
  input clk;
  input arst_n;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for bbox_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg  state_var;
  reg  state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : bbox_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_staller
// ------------------------------------------------------------------


module bbox_core_staller (
  clk, arst_n, core_wen, core_wten, bbox_req_stream_rsci_wen_comp, bbox_resp_stream_rsci_wen_comp,
      core_flen_unreg
);
  input clk;
  input arst_n;
  output core_wen;
  output core_wten;
  input bbox_req_stream_rsci_wen_comp;
  input bbox_resp_stream_rsci_wen_comp;
  input core_flen_unreg;


  // Interconnect Declarations
  reg core_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign core_wen = bbox_req_stream_rsci_wen_comp & bbox_resp_stream_rsci_wen_comp
      & (~ core_flen_unreg);
  assign core_wten = core_wten_reg;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      core_wten_reg <= 1'b0;
    end
    else begin
      core_wten_reg <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_23_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_23
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_23_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_23
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_23_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_23_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_23_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_23_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_23_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_23_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_23_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_23_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_23_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_23_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_23_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_23_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_23_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_23_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_23_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_23_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_23_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_23_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_23_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_23_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_23
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_23_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_23
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_23_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_23_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_23_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_23_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_23_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_23_cs_lp_piped_fp_mult_23_8_0_cmp_23_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_23_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_23_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_23_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_23_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_23_cs_lp_piped_fp_mult_23_8_0_cmp_23_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_23_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_23_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_cs_lp_piped_fp_mult_23_8_0_cmp_23_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_cs_lp_piped_fp_mult_23_8_0_cmp_23_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_23_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_23_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_23_cs_lp_piped_fp_mult_23_8_0_cmp_23_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_23_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_23_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_22
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_22
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_22_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_22_a_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_b_core, ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_22_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_a, ccs_lp_piped_fp_mult_23_8_0_cmp_22_b,
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_22_bawt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_22_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_22_bdwt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_a;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_b;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_22_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_22_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_22_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_22_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_22_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_bcwt);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_22_a = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_22_a_core[30:16])
      , 16'b0000000000000000};
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_22_b = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_22_b_core[30:23])
      , 23'b00000000000000000000000};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_22_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_22_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_22_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_22_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_22_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_22_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_22_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_22
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_22
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_22_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_22_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_22_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_22_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_22_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_22_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_22_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_22_cs_lp_piped_fp_mult_23_8_0_cmp_22_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_22_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_22_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_22_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_22_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_22_cs_lp_piped_fp_mult_23_8_0_cmp_22_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_22_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_22_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_cs_lp_piped_fp_mult_23_8_0_cmp_22_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_cs_lp_piped_fp_mult_23_8_0_cmp_22_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_22_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_22_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_22_cs_lp_piped_fp_mult_23_8_0_cmp_22_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_22_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_22_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_21_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_21
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_21_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_21
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_21_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_21_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_21_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_21_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_21_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_21_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_21_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_21_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_3_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_3_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_21_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_21_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_21_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_21_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_21_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_21_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_21_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_3_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_21_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_21_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_3_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_3_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_21_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_3_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_21_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_21_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_21
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_21_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_21
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_21_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_21_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_21_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_21_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_21_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_21_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_21_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_21_cs_lp_piped_fp_mult_23_8_0_cmp_21_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_21_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_21_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_3_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_3_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_21_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_21_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_21_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_21_cs_lp_piped_fp_mult_23_8_0_cmp_21_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_21_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_21_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_cs_lp_piped_fp_mult_23_8_0_cmp_21_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_cs_lp_piped_fp_mult_23_8_0_cmp_21_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_21_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_3_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_21_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_21_cs_lp_piped_fp_mult_23_8_0_cmp_21_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_3_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_3_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_21_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_3_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_21_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_20
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_20
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_20_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_20_a_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_b_core, ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_20_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_a, ccs_lp_piped_fp_mult_23_8_0_cmp_20_b,
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_20_bawt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_20_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_20_bdwt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_a;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_b;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_20_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_4_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_4_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_20_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_20_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_20_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_20_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_bcwt);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_20_a = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_20_a_core[30:16])
      , 16'b0000000000000000};
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_20_b = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_20_b_core[30:23])
      , 23'b00000000000000000000000};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_20_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_20_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_20_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_4_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_20_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_20_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_4_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_4_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_20_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_4_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_20_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_20
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_20
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_20_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_20_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_20_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_20_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_20_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_20_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_20_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_20_cs_lp_piped_fp_mult_23_8_0_cmp_20_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_20_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_4_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_4_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_20_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_20_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_20_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_20_cs_lp_piped_fp_mult_23_8_0_cmp_20_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_20_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_20_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_cs_lp_piped_fp_mult_23_8_0_cmp_20_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_cs_lp_piped_fp_mult_23_8_0_cmp_20_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_20_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_4_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_20_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_20_cs_lp_piped_fp_mult_23_8_0_cmp_20_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_4_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_4_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_20_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_4_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_20_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_19_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_19
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_19_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_19
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_19_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_19_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_19_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_19_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_19_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_19_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_19_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_19_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_5_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_5_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_19_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_19_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_19_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_19_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_19_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_19_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_19_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_5_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_19_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_19_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_5_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_5_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_19_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_5_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_19_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_19_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_19
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_19_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_19
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_19_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_19_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_19_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_19_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_19_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_19_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_19_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_19_cs_lp_piped_fp_mult_23_8_0_cmp_19_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_19_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_19_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_5_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_5_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_19_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_19_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_19_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_19_cs_lp_piped_fp_mult_23_8_0_cmp_19_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_19_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_19_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_cs_lp_piped_fp_mult_23_8_0_cmp_19_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_cs_lp_piped_fp_mult_23_8_0_cmp_19_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_19_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_5_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_19_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_19_cs_lp_piped_fp_mult_23_8_0_cmp_19_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_5_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_5_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_19_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_5_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_19_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_18
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_18
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_18_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_18_a_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_b_core, ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_18_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_a, ccs_lp_piped_fp_mult_23_8_0_cmp_18_b,
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_18_bawt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_18_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_18_bdwt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_a;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_b;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_18_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_6_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_6_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_18_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_18_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_18_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_18_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_bcwt);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_18_a = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_18_a_core[30:16])
      , 16'b0000000000000000};
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_18_b = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_18_b_core[30:23])
      , 23'b00000000000000000000000};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_18_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_18_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_18_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_6_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_18_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_18_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_6_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_6_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_18_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_6_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_18_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_18
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_18
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_18_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_18_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_18_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_18_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_18_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_18_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_18_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_18_cs_lp_piped_fp_mult_23_8_0_cmp_18_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_18_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_6_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_6_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_18_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_18_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_18_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_18_cs_lp_piped_fp_mult_23_8_0_cmp_18_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_18_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_18_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_cs_lp_piped_fp_mult_23_8_0_cmp_18_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_cs_lp_piped_fp_mult_23_8_0_cmp_18_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_18_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_6_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_18_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_18_cs_lp_piped_fp_mult_23_8_0_cmp_18_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_6_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_6_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_18_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_6_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_18_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_17_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_17
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_17_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_17
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_17_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_17_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_17_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_17_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_17_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_17_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_17_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_17_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_7_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_7_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_17_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_17_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_17_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_17_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_17_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_17_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_17_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_7_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_17_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_17_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_7_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_7_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_17_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_7_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_17_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_17_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_17
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_17_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_17
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_17_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_17_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_17_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_17_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_17_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_17_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_17_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_17_cs_lp_piped_fp_mult_23_8_0_cmp_17_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_17_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_17_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_7_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_7_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_17_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_17_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_17_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_17_cs_lp_piped_fp_mult_23_8_0_cmp_17_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_17_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_17_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_cs_lp_piped_fp_mult_23_8_0_cmp_17_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_cs_lp_piped_fp_mult_23_8_0_cmp_17_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_17_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_7_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_17_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_17_cs_lp_piped_fp_mult_23_8_0_cmp_17_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_7_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_7_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_17_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_7_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_17_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_16
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_16
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_16_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_16_a_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_b_core, ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_16_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_a, ccs_lp_piped_fp_mult_23_8_0_cmp_16_b,
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_16_bawt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_16_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_16_bdwt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_a;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_b;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_16_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_8_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_8_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_16_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_16_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_16_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_16_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_bcwt);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_16_a = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_16_a_core[30:16])
      , 16'b0000000000000000};
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_16_b = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_16_b_core[30:23])
      , 23'b00000000000000000000000};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_16_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_16_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_16_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_8_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_16_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_16_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_8_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_8_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_16_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_8_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_16_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_16
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_16
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_16_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_16_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_16_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_16_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_16_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_16_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_16_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_16_cs_lp_piped_fp_mult_23_8_0_cmp_16_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_16_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_8_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_8_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_16_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_16_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_16_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_16_cs_lp_piped_fp_mult_23_8_0_cmp_16_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_16_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_16_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_cs_lp_piped_fp_mult_23_8_0_cmp_16_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_cs_lp_piped_fp_mult_23_8_0_cmp_16_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_16_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_8_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_16_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_16_cs_lp_piped_fp_mult_23_8_0_cmp_16_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_8_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_8_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_16_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_8_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_16_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_15_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_15
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_15_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_15
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_15_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_15_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_15_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_15_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_15_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_15_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_15_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_15_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_9_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_9_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_15_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_15_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_15_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_15_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_15_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_15_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_15_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_9_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_15_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_15_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_9_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_9_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_15_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_9_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_15_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_15_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_15
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_15_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_15
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_15_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_15_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_15_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_15_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_15_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_15_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_15_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_15_cs_lp_piped_fp_mult_23_8_0_cmp_15_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_15_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_15_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_9_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_9_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_15_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_15_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_15_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_15_cs_lp_piped_fp_mult_23_8_0_cmp_15_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_15_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_15_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_cs_lp_piped_fp_mult_23_8_0_cmp_15_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_cs_lp_piped_fp_mult_23_8_0_cmp_15_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_15_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_9_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_15_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_15_cs_lp_piped_fp_mult_23_8_0_cmp_15_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_9_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_9_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_15_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_9_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_15_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_14
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_14
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_14_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_14_a_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_b_core, ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_14_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_a, ccs_lp_piped_fp_mult_23_8_0_cmp_14_b,
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_14_bawt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_14_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_14_bdwt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_a;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_b;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_14_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_10_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_10_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_14_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_14_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_14_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_14_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_bcwt);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_14_a = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_14_a_core[30:16])
      , 16'b0000000000000000};
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_14_b = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_14_b_core[30:23])
      , 23'b00000000000000000000000};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_14_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_14_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_14_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_10_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_14_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_14_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_10_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_10_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_14_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_10_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_14_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_14
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_14
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_14_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_14_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_14_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_14_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_14_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_14_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_14_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_14_cs_lp_piped_fp_mult_23_8_0_cmp_14_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_14_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_10_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_10_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_14_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_14_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_14_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_14_cs_lp_piped_fp_mult_23_8_0_cmp_14_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_14_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_14_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_cs_lp_piped_fp_mult_23_8_0_cmp_14_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_cs_lp_piped_fp_mult_23_8_0_cmp_14_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_14_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_10_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_14_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_14_cs_lp_piped_fp_mult_23_8_0_cmp_14_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_10_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_10_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_14_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_10_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_14_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_13_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_13
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_13_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_13
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_13_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_13_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_13_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_13_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_13_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_13_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_13_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_13_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_11_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_11_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_13_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_13_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_13_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_13_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_13_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_13_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_13_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_11_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_13_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_13_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_11_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_11_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_13_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_11_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_13_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_13_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_13
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_13_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_13
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_13_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_13_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_13_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_13_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_13_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_13_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_13_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_13_cs_lp_piped_fp_mult_23_8_0_cmp_13_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_13_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_13_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_11_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_11_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_13_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_13_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_13_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_13_cs_lp_piped_fp_mult_23_8_0_cmp_13_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_13_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_13_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_cs_lp_piped_fp_mult_23_8_0_cmp_13_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_cs_lp_piped_fp_mult_23_8_0_cmp_13_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_13_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_11_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_13_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_13_cs_lp_piped_fp_mult_23_8_0_cmp_13_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_11_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_11_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_13_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_11_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_13_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_12
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_12
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_12_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_12_a_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_b_core, ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_12_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_a, ccs_lp_piped_fp_mult_23_8_0_cmp_12_b,
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_12_bawt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_12_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_12_bdwt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_a;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_b;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_12_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_12_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_12_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_12_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_12_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_12_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_12_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_bcwt);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_12_a = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_12_a_core[30:16])
      , 16'b0000000000000000};
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_12_b = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_12_b_core[30:23])
      , 23'b00000000000000000000000};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_12_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_12_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_12_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_12_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_12_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_12_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_12_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_12_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_12_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_12_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_12_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_12
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_12
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_12_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_12_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_12_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_12_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_12_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_12_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_12_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_12_cs_lp_piped_fp_mult_23_8_0_cmp_12_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_12_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_12_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_12_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_12_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_12_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_12_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_12_cs_lp_piped_fp_mult_23_8_0_cmp_12_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_12_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_12_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_cs_lp_piped_fp_mult_23_8_0_cmp_12_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_cs_lp_piped_fp_mult_23_8_0_cmp_12_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_12_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_12_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_12_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_12_cs_lp_piped_fp_mult_23_8_0_cmp_12_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_12_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_12_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_12_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_12_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_12_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_11_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_11
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_11_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_11
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_11_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_11_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_11_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_11_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_11_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_11_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_11_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_11_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_13_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_13_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_11_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_11_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_11_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_11_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_11_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_11_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_11_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_13_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_11_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_11_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_13_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_13_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_11_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_13_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_11_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_11_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_11
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_11_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_11
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_11_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_11_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_11_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_11_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_11_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_11_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_11_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_11_cs_lp_piped_fp_mult_23_8_0_cmp_11_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_11_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_11_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_13_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_13_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_11_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_11_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_11_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_11_cs_lp_piped_fp_mult_23_8_0_cmp_11_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_11_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_11_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_cs_lp_piped_fp_mult_23_8_0_cmp_11_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_cs_lp_piped_fp_mult_23_8_0_cmp_11_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_11_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_13_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_11_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_11_cs_lp_piped_fp_mult_23_8_0_cmp_11_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_13_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_13_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_11_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_13_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_11_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_10
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_10
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_10_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_10_a_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_b_core, ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_10_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_a, ccs_lp_piped_fp_mult_23_8_0_cmp_10_b,
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_10_bawt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_10_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_10_bdwt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_a;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_b;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_10_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_14_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_14_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_10_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_10_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_10_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_10_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_bcwt);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_10_a = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_10_a_core[30:16])
      , 16'b0000000000000000};
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_10_b = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_10_b_core[30:23])
      , 23'b00000000000000000000000};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_10_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_10_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_10_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_14_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_10_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_10_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_14_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_14_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_10_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_14_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_10_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_10
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_10
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_10_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_10_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_10_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_10_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_10_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_10_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_10_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_10_cs_lp_piped_fp_mult_23_8_0_cmp_10_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_10_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_14_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_14_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_10_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_10_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_10_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_10_cs_lp_piped_fp_mult_23_8_0_cmp_10_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_10_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_10_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_cs_lp_piped_fp_mult_23_8_0_cmp_10_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_cs_lp_piped_fp_mult_23_8_0_cmp_10_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_10_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_14_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_10_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_10_cs_lp_piped_fp_mult_23_8_0_cmp_10_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_14_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_14_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_10_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_14_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_10_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_9_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_9
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_9_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_9
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_9_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_9_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_9_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_9_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_9_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_9_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_9_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_9_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_15_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_15_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_9_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_9_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_9_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_9_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_9_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_9_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_9_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_15_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_9_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_9_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_15_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_15_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_9_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_15_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_9_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_9_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_9
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_9_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_9
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_9_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_9_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_9_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_9_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_9_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_9_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_9_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_9_cs_lp_piped_fp_mult_23_8_0_cmp_9_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_9_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_9_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_15_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_15_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_9_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_9_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_9_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_9_cs_lp_piped_fp_mult_23_8_0_cmp_9_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_9_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_9_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_cs_lp_piped_fp_mult_23_8_0_cmp_9_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_cs_lp_piped_fp_mult_23_8_0_cmp_9_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_9_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_15_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_9_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_9_cs_lp_piped_fp_mult_23_8_0_cmp_9_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_15_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_15_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_9_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_15_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_9_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_8
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_8
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_8_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_8_a_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_b_core, ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_8_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_a, ccs_lp_piped_fp_mult_23_8_0_cmp_8_b, ccs_lp_piped_fp_mult_23_8_0_cmp_8_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_8_bawt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_8_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_8_bdwt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_a;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_b;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_8_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_16_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_16_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_8_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_8_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_8_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_8_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_bcwt);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_8_a = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_8_a_core[30:16])
      , 16'b0000000000000000};
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_8_b = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_8_b_core[30:23])
      , 23'b00000000000000000000000};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_8_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_8_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_8_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_16_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_8_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_8_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_16_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_16_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_8_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_16_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_8_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_8
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_8
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_8_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_8_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_8_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_8_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_8_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_8_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_8_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_8_cs_lp_piped_fp_mult_23_8_0_cmp_8_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_8_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_16_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_16_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_8_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_8_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_8_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_8_cs_lp_piped_fp_mult_23_8_0_cmp_8_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_8_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_8_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_cs_lp_piped_fp_mult_23_8_0_cmp_8_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_cs_lp_piped_fp_mult_23_8_0_cmp_8_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_8_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_16_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_8_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_8_cs_lp_piped_fp_mult_23_8_0_cmp_8_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_16_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_16_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_8_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_16_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_8_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_7_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_7
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_7_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_7
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_7_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_7_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_7_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_7_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_7_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_7_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_7_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_7_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_17_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_17_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_7_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_7_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_7_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_7_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_7_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_7_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_7_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_17_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_7_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_7_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_17_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_17_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_7_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_17_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_7_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_7_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_7
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_7_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_7
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_7_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_7_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_7_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_7_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_7_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_7_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_7_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_7_cs_lp_piped_fp_mult_23_8_0_cmp_7_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_7_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_7_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_17_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_17_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_7_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_7_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_7_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_7_cs_lp_piped_fp_mult_23_8_0_cmp_7_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_7_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_7_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_cs_lp_piped_fp_mult_23_8_0_cmp_7_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_cs_lp_piped_fp_mult_23_8_0_cmp_7_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_7_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_17_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_7_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_7_cs_lp_piped_fp_mult_23_8_0_cmp_7_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_17_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_17_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_7_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_17_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_7_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_6
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_6
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_6_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_6_a_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_b_core, ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_6_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_a, ccs_lp_piped_fp_mult_23_8_0_cmp_6_b, ccs_lp_piped_fp_mult_23_8_0_cmp_6_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_6_bawt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_6_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_6_bdwt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_a;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_b;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_6_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_18_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_18_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_6_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_6_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_6_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_6_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_bcwt);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_6_a = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_6_a_core[30:16])
      , 16'b0000000000000000};
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_6_b = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_6_b_core[30:23])
      , 23'b00000000000000000000000};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_6_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_6_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_6_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_18_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_6_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_6_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_18_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_18_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_6_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_18_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_6_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_6
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_6
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_6_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_6_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_6_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_6_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_6_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_6_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_6_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_6_cs_lp_piped_fp_mult_23_8_0_cmp_6_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_6_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_18_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_18_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_6_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_6_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_6_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_6_cs_lp_piped_fp_mult_23_8_0_cmp_6_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_6_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_6_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_cs_lp_piped_fp_mult_23_8_0_cmp_6_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_cs_lp_piped_fp_mult_23_8_0_cmp_6_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_6_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_18_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_6_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_6_cs_lp_piped_fp_mult_23_8_0_cmp_6_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_18_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_18_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_6_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_18_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_6_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_5
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_5
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_5_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_5_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_5_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_5_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_5_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_5_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_5_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_5_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_19_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_19_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_5_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_5_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_5_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_5_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_5_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_5_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_5_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_19_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_5_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_5_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_19_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_19_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_5_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_19_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_5_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_5
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_5
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_5_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_5_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_5_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_5_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_5_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_5_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_5_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_5_cs_lp_piped_fp_mult_23_8_0_cmp_5_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_5_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_5_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_19_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_19_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_5_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_5_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_5_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_5_cs_lp_piped_fp_mult_23_8_0_cmp_5_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_5_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_5_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_cs_lp_piped_fp_mult_23_8_0_cmp_5_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_cs_lp_piped_fp_mult_23_8_0_cmp_5_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_5_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_19_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_5_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_5_cs_lp_piped_fp_mult_23_8_0_cmp_5_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_19_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_19_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_5_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_19_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_5_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_4
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_4
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_4_a_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_b_core, ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_4_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_a, ccs_lp_piped_fp_mult_23_8_0_cmp_4_b, ccs_lp_piped_fp_mult_23_8_0_cmp_4_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_4_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_4_bdwt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_a;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_b;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_4_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_20_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_20_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_4_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_4_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_4_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_bcwt);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_4_a = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_4_a_core[30:16])
      , 16'b0000000000000000};
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_4_b = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_4_b_core[30:23])
      , 23'b00000000000000000000000};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_4_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_4_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_4_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_20_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_4_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_4_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_20_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_20_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_4_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_20_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_4_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_4
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_4
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_4_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_4_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_4_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_4_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_4_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_4_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_4_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_4_cs_lp_piped_fp_mult_23_8_0_cmp_4_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_4_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_20_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_20_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_4_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_4_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_4_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_4_cs_lp_piped_fp_mult_23_8_0_cmp_4_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_4_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_4_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_cs_lp_piped_fp_mult_23_8_0_cmp_4_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_cs_lp_piped_fp_mult_23_8_0_cmp_4_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_4_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_20_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_4_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_4_cs_lp_piped_fp_mult_23_8_0_cmp_4_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_20_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_20_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_4_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_20_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_4_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_3_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_3
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_3_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_3
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_3_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_3_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_3_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_3_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_3_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_3_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_3_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_3_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_21_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_21_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_3_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_3_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_3_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_3_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_3_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_3_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_3_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_21_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_3_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_3_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_21_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_21_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_3_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_21_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_3_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_3_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_3
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_3_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_3
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_3_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_3_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_3_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_3_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_3_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_3_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_3_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_3_cs_lp_piped_fp_mult_23_8_0_cmp_3_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_3_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_3_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_21_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_21_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_3_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_3_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_3_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_3_cs_lp_piped_fp_mult_23_8_0_cmp_3_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_3_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_3_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_cs_lp_piped_fp_mult_23_8_0_cmp_3_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_cs_lp_piped_fp_mult_23_8_0_cmp_3_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_3_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_21_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_3_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_3_cs_lp_piped_fp_mult_23_8_0_cmp_3_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_21_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_21_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_3_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_21_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_3_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_2
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_2
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_2_a_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_b_core, ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_a, ccs_lp_piped_fp_mult_23_8_0_cmp_2_b, ccs_lp_piped_fp_mult_23_8_0_cmp_2_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_a;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_b;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_2_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_22_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_22_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_2_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_2_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_bcwt);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_2_a = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_2_a_core[30:16])
      , 16'b0000000000000000};
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_2_b = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_2_b_core[30:23])
      , 23'b00000000000000000000000};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_2_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_2_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_22_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_22_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_22_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_2_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_22_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_2_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_2
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_2
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_2_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_2_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_2_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_2_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_2_cs_lp_piped_fp_mult_23_8_0_cmp_2_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_2_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_22_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_22_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_2_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_2_cs_lp_piped_fp_mult_23_8_0_cmp_2_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_2_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_2_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_cs_lp_piped_fp_mult_23_8_0_cmp_2_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_cs_lp_piped_fp_mult_23_8_0_cmp_2_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_2_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_22_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_2_cs_lp_piped_fp_mult_23_8_0_cmp_2_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_22_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_22_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_2_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_22_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_2_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_1
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_1
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_1_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_23_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_23_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_1_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_1_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_1_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_1_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_23_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_23_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_23_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_1_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_23_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_1_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_1
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_1
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_1_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_1_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_1_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_1_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_1_cs_lp_piped_fp_mult_23_8_0_cmp_1_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_1_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_23_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_23_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_1_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_1_cs_lp_piped_fp_mult_23_8_0_cmp_1_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_1_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_1_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_cs_lp_piped_fp_mult_23_8_0_cmp_1_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_cs_lp_piped_fp_mult_23_8_0_cmp_1_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_1_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_23_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_1_cs_lp_piped_fp_mult_23_8_0_cmp_1_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_23_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_23_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_1_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_23_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_1_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_a_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_b_core, ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_a, ccs_lp_piped_fp_mult_23_8_0_cmp_b, ccs_lp_piped_fp_mult_23_8_0_cmp_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_bawt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_a;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_b;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_bcwt);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_a = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_a_core[30:16])
      , 16'b0000000000000000};
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_b = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_b_core[30:23])
      , 23'b00000000000000000000000};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_oswt_unreg, ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_launch_core_sct, ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_cs_lp_piped_fp_mult_23_8_0_cmp_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_cs_lp_piped_fp_mult_23_8_0_cmp_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_cs_lp_piped_fp_mult_23_8_0_cmp_pdswt0 <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_cs_lp_piped_fp_mult_23_8_0_cmp_pdswt0 <= (~
          core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_cs_lp_piped_fp_mult_23_8_0_cmp_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_11_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_11
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_11_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_11
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_11_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_11_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_11_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_11_bdwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_11_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_11_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_11_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_11_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_11_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_11_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_11_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_11_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_11_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_11_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_11_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_11_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_11_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_11_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_11_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_11_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_11_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_11_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_11_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_11_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_11_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_11_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_11_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_11_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_11_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_11_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_11_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_11_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_11_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_11_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_11_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_11_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_11_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_11
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_11_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_11
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_11_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_11_biwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_11_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_11_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_11_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_11_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_11_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_11_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_11_cs_lp_piped_fp_add_23_8_0_cmp_11_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_11_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_11_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_11_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_11_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_11_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_11_cs_lp_piped_fp_add_23_8_0_cmp_11_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_11_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_11_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_11_cs_lp_piped_fp_add_23_8_0_cmp_11_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_11_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_11_cs_lp_piped_fp_add_23_8_0_cmp_11_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_11_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_11_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_11_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_11_cs_lp_piped_fp_add_23_8_0_cmp_11_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_11_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_11_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_10_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_10
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_10_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_10
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_10_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_10_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_10_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_10_bdwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_10_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_10_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_10_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_10_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_10_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_10_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_10_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_10_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_10_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_10_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_10_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_10_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_10_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_10_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_10_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_10_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_10_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_10_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_10_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_10_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_10_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_10_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_10_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_10_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_10_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_10_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_10_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_10_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_10_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_10_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_10_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_10_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_10_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_10
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_10_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_10
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_10_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_10_biwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_10_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_10_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_10_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_10_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_10_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_10_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_10_cs_lp_piped_fp_add_23_8_0_cmp_10_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_10_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_10_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_10_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_10_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_10_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_10_cs_lp_piped_fp_add_23_8_0_cmp_10_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_10_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_10_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_10_cs_lp_piped_fp_add_23_8_0_cmp_10_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_10_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_10_cs_lp_piped_fp_add_23_8_0_cmp_10_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_10_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_10_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_10_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_10_cs_lp_piped_fp_add_23_8_0_cmp_10_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_10_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_10_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_9_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_9
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_9_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_9
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_9_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_9_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_9_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_9_bdwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_9_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_9_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_9_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_9_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_9_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_9_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_9_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_9_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_9_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_9_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_3_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_3_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_9_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_9_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_9_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_9_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_9_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_9_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_9_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_9_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_9_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_9_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_9_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_9_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_9_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_9_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_9_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_9_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_9_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_9_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_3_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_9_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_9_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_3_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_3_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_9_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_3_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_9_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_9_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_9
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_9_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_9
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_9_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_9_biwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_9_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_9_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_9_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_9_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_9_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_9_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_9_cs_lp_piped_fp_add_23_8_0_cmp_9_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_9_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_9_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_3_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_3_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_9_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_9_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_9_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_9_cs_lp_piped_fp_add_23_8_0_cmp_9_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_9_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_9_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_9_cs_lp_piped_fp_add_23_8_0_cmp_9_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_9_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_9_cs_lp_piped_fp_add_23_8_0_cmp_9_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_9_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_9_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_3_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_9_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_9_cs_lp_piped_fp_add_23_8_0_cmp_9_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_3_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_3_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_9_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_3_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_9_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_8_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_8
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_8_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_8
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_8_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_8_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_8_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_8_bdwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_8_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_8_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_8_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_8_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_8_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_8_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_8_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_8_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_8_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_8_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_4_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_4_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_8_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_8_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_8_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_8_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_8_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_8_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_8_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_8_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_8_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_8_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_8_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_8_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_8_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_8_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_8_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_8_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_8_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_8_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_4_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_8_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_8_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_4_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_4_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_8_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_4_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_8_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_8_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_8
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_8_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_8
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_8_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_8_biwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_8_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_8_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_8_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_8_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_8_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_8_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_8_cs_lp_piped_fp_add_23_8_0_cmp_8_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_8_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_8_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_4_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_4_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_8_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_8_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_8_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_8_cs_lp_piped_fp_add_23_8_0_cmp_8_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_8_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_8_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_8_cs_lp_piped_fp_add_23_8_0_cmp_8_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_8_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_8_cs_lp_piped_fp_add_23_8_0_cmp_8_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_8_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_8_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_4_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_8_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_8_cs_lp_piped_fp_add_23_8_0_cmp_8_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_4_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_4_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_8_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_4_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_8_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_7_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_7
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_7_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_7
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_7_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_7_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_7_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_7_bdwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_7_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_7_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_7_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_7_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_7_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_7_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_7_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_7_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_7_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_7_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_5_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_5_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_7_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_7_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_7_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_7_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_7_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_7_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_7_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_7_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_7_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_7_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_7_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_7_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_7_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_7_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_7_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_7_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_7_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_7_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_5_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_7_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_7_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_5_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_5_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_7_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_5_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_7_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_7_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_7
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_7_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_7
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_7_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_7_biwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_7_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_7_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_7_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_7_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_7_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_7_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_7_cs_lp_piped_fp_add_23_8_0_cmp_7_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_7_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_7_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_5_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_5_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_7_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_7_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_7_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_7_cs_lp_piped_fp_add_23_8_0_cmp_7_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_7_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_7_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_7_cs_lp_piped_fp_add_23_8_0_cmp_7_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_7_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_7_cs_lp_piped_fp_add_23_8_0_cmp_7_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_7_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_7_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_5_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_7_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_7_cs_lp_piped_fp_add_23_8_0_cmp_7_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_5_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_5_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_7_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_5_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_7_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_6_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_6
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_6_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_6
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_6_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_6_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_6_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_6_bdwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_6_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_6_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_6_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_6_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_6_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_6_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_6_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_6_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_6_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_6_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_6_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_6_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_6_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_6_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_6_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_6_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_6_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_6_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_6_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_6_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_6_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_6_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_6_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_6_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_6_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_6_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_6_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_6_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_6_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_6_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_6_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_6_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_6_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_6_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_6_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_6_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_6_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_6_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_6_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_6
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_6_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_6
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_6_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_6_biwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_6_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_6_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_6_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_6_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_6_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_6_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_6_cs_lp_piped_fp_add_23_8_0_cmp_6_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_6_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_6_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_6_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_6_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_6_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_6_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_6_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_6_cs_lp_piped_fp_add_23_8_0_cmp_6_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_6_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_6_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_6_cs_lp_piped_fp_add_23_8_0_cmp_6_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_6_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_6_cs_lp_piped_fp_add_23_8_0_cmp_6_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_6_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_6_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_6_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_6_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_6_cs_lp_piped_fp_add_23_8_0_cmp_6_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_6_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_6_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_6_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_6_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_6_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_5_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_5
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_5_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_5
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_5_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_5_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_5_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_5_bdwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_5_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_5_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_5_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_5_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_5_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_5_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_5_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_5_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_5_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_5_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_7_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_7_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_5_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_5_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_5_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_5_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_5_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_5_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_5_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_5_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_5_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_5_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_5_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_5_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_5_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_5_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_5_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_5_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_5_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_5_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_7_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_5_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_5_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_7_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_7_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_5_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_7_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_5_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_5_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_5
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_5_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_5
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_5_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_5_biwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_5_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_5_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_5_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_5_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_5_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_5_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_5_cs_lp_piped_fp_add_23_8_0_cmp_5_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_5_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_5_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_7_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_7_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_5_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_5_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_5_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_5_cs_lp_piped_fp_add_23_8_0_cmp_5_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_5_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_5_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_5_cs_lp_piped_fp_add_23_8_0_cmp_5_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_5_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_5_cs_lp_piped_fp_add_23_8_0_cmp_5_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_5_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_5_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_7_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_5_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_5_cs_lp_piped_fp_add_23_8_0_cmp_5_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_7_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_7_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_5_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_7_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_5_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_4_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_4
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_4_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_4
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_4_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_4_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_4_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_4_bdwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_4_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_4_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_4_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_4_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_4_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_4_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_4_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_4_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_4_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_4_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_8_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_8_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_4_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_4_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_4_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_4_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_4_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_4_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_4_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_4_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_4_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_4_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_4_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_4_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_4_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_4_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_4_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_4_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_4_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_4_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_8_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_4_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_4_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_8_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_8_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_4_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_8_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_4_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_4_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_4
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_4_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_4
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_4_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_4_biwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_4_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_4_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_4_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_4_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_4_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_4_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_4_cs_lp_piped_fp_add_23_8_0_cmp_4_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_4_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_4_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_8_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_8_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_4_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_4_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_4_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_4_cs_lp_piped_fp_add_23_8_0_cmp_4_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_4_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_4_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_4_cs_lp_piped_fp_add_23_8_0_cmp_4_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_4_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_4_cs_lp_piped_fp_add_23_8_0_cmp_4_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_4_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_4_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_8_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_4_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_4_cs_lp_piped_fp_add_23_8_0_cmp_4_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_8_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_8_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_4_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_8_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_4_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_3_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_3
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_3_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_3
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_3_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_3_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_3_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_3_bdwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_3_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_3_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_3_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_3_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_3_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_3_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_3_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_3_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_3_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_3_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_9_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_9_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_3_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_3_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_3_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_3_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_3_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_3_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_3_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_3_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_3_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_3_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_3_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_3_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_3_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_3_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_3_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_3_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_3_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_3_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_9_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_3_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_3_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_9_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_9_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_3_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_9_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_3_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_3_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_3
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_3_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_3
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_3_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_3_biwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_3_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_3_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_3_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_3_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_3_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_3_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_3_cs_lp_piped_fp_add_23_8_0_cmp_3_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_3_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_3_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_9_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_9_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_3_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_3_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_3_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_3_cs_lp_piped_fp_add_23_8_0_cmp_3_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_3_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_3_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_3_cs_lp_piped_fp_add_23_8_0_cmp_3_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_3_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_3_cs_lp_piped_fp_add_23_8_0_cmp_3_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_3_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_3_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_9_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_3_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_3_cs_lp_piped_fp_add_23_8_0_cmp_3_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_9_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_9_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_3_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_9_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_3_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_2
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_2
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_2_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_2_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_10_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_10_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_2_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_2_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_2_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_2_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_2_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_2_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_2_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_2_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_2_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_2_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_2_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_2_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_2_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_2_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_10_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_10_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_10_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_2_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_10_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_2_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_2
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_2
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_2_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_2_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_2_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_2_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_2_cs_lp_piped_fp_add_23_8_0_cmp_2_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_2_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_10_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_10_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_2_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_2_cs_lp_piped_fp_add_23_8_0_cmp_2_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_2_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_2_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_2_cs_lp_piped_fp_add_23_8_0_cmp_2_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_2_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_2_cs_lp_piped_fp_add_23_8_0_cmp_2_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_2_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_2_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_10_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_2_cs_lp_piped_fp_add_23_8_0_cmp_2_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_10_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_10_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_2_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_10_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_2_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_1
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_1
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_1_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_1_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_11_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_11_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_1_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_1_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_1_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_1_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_1_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_1_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_1_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_1_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_1_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_1_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_1_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_1_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_1_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_1_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_11_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_11_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_11_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_1_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_11_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_1_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_1
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_1
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_1_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_1_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_1_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_1_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_1_cs_lp_piped_fp_add_23_8_0_cmp_1_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_1_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_11_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_11_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_1_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_1_cs_lp_piped_fp_add_23_8_0_cmp_1_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_1_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_1_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_1_cs_lp_piped_fp_add_23_8_0_cmp_1_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_1_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_1_cs_lp_piped_fp_add_23_8_0_cmp_1_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_1_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_1_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_11_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_1_cs_lp_piped_fp_add_23_8_0_cmp_1_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_11_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_11_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_1_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_11_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_1_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_oswt_unreg, ccs_lp_piped_fp_add_23_8_0_cmp_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_cs_lp_piped_fp_add_23_8_0_cmp_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_cs_lp_piped_fp_add_23_8_0_cmp_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_cs_lp_piped_fp_add_23_8_0_cmp_pdswt0 <= 1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_cs_lp_piped_fp_add_23_8_0_cmp_pdswt0 <= (~ core_wten)
          & ccs_lp_piped_fp_add_23_8_0_cmp_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_cs_lp_piped_fp_add_23_8_0_cmp_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_bbox_resp_stream_rsci_bbox_resp_stream_wait_dp
// ------------------------------------------------------------------


module bbox_core_bbox_resp_stream_rsci_bbox_resp_stream_wait_dp (
  clk, arst_n, bbox_resp_stream_rsci_oswt_unreg, bbox_resp_stream_rsci_bawt, bbox_resp_stream_rsci_wen_comp,
      bbox_resp_stream_rsci_biwt, bbox_resp_stream_rsci_bdwt, bbox_resp_stream_rsci_bcwt
);
  input clk;
  input arst_n;
  input bbox_resp_stream_rsci_oswt_unreg;
  output bbox_resp_stream_rsci_bawt;
  output bbox_resp_stream_rsci_wen_comp;
  input bbox_resp_stream_rsci_biwt;
  input bbox_resp_stream_rsci_bdwt;
  output bbox_resp_stream_rsci_bcwt;
  reg bbox_resp_stream_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign bbox_resp_stream_rsci_bawt = bbox_resp_stream_rsci_biwt | bbox_resp_stream_rsci_bcwt;
  assign bbox_resp_stream_rsci_wen_comp = (~ bbox_resp_stream_rsci_oswt_unreg) |
      bbox_resp_stream_rsci_bawt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      bbox_resp_stream_rsci_bcwt <= 1'b0;
    end
    else begin
      bbox_resp_stream_rsci_bcwt <= ~((~(bbox_resp_stream_rsci_bcwt | bbox_resp_stream_rsci_biwt))
          | bbox_resp_stream_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_bbox_resp_stream_rsci_bbox_resp_stream_wait_ctrl
// ------------------------------------------------------------------


module bbox_core_bbox_resp_stream_rsci_bbox_resp_stream_wait_ctrl (
  core_wen, bbox_resp_stream_rsci_oswt_unreg, bbox_resp_stream_rsci_iswt0, bbox_resp_stream_rsci_biwt,
      bbox_resp_stream_rsci_bdwt, bbox_resp_stream_rsci_bcwt, bbox_resp_stream_rsci_irdy,
      bbox_resp_stream_rsci_ivld_core_sct
);
  input core_wen;
  input bbox_resp_stream_rsci_oswt_unreg;
  input bbox_resp_stream_rsci_iswt0;
  output bbox_resp_stream_rsci_biwt;
  output bbox_resp_stream_rsci_bdwt;
  input bbox_resp_stream_rsci_bcwt;
  input bbox_resp_stream_rsci_irdy;
  output bbox_resp_stream_rsci_ivld_core_sct;


  // Interconnect Declarations
  wire bbox_resp_stream_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign bbox_resp_stream_rsci_bdwt = bbox_resp_stream_rsci_oswt_unreg & core_wen;
  assign bbox_resp_stream_rsci_biwt = bbox_resp_stream_rsci_ogwt & bbox_resp_stream_rsci_irdy;
  assign bbox_resp_stream_rsci_ogwt = bbox_resp_stream_rsci_iswt0 & (~ bbox_resp_stream_rsci_bcwt);
  assign bbox_resp_stream_rsci_ivld_core_sct = bbox_resp_stream_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_bbox_req_stream_rsci_bbox_req_stream_wait_dp
// ------------------------------------------------------------------


module bbox_core_bbox_req_stream_rsci_bbox_req_stream_wait_dp (
  clk, arst_n, bbox_req_stream_rsci_oswt_unreg, bbox_req_stream_rsci_bawt, bbox_req_stream_rsci_wen_comp,
      bbox_req_stream_rsci_idat_mxwt, bbox_req_stream_rsci_biwt, bbox_req_stream_rsci_bdwt,
      bbox_req_stream_rsci_bcwt, bbox_req_stream_rsci_idat
);
  input clk;
  input arst_n;
  input bbox_req_stream_rsci_oswt_unreg;
  output bbox_req_stream_rsci_bawt;
  output bbox_req_stream_rsci_wen_comp;
  output [385:0] bbox_req_stream_rsci_idat_mxwt;
  input bbox_req_stream_rsci_biwt;
  input bbox_req_stream_rsci_bdwt;
  output bbox_req_stream_rsci_bcwt;
  reg bbox_req_stream_rsci_bcwt;
  input [385:0] bbox_req_stream_rsci_idat;


  // Interconnect Declarations
  reg [385:0] bbox_req_stream_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign bbox_req_stream_rsci_bawt = bbox_req_stream_rsci_biwt | bbox_req_stream_rsci_bcwt;
  assign bbox_req_stream_rsci_wen_comp = (~ bbox_req_stream_rsci_oswt_unreg) | bbox_req_stream_rsci_bawt;
  assign bbox_req_stream_rsci_idat_mxwt = MUX_v_386_2_2(bbox_req_stream_rsci_idat,
      bbox_req_stream_rsci_idat_bfwt, bbox_req_stream_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      bbox_req_stream_rsci_bcwt <= 1'b0;
    end
    else begin
      bbox_req_stream_rsci_bcwt <= ~((~(bbox_req_stream_rsci_bcwt | bbox_req_stream_rsci_biwt))
          | bbox_req_stream_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      bbox_req_stream_rsci_idat_bfwt <= 386'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( bbox_req_stream_rsci_biwt ) begin
      bbox_req_stream_rsci_idat_bfwt <= bbox_req_stream_rsci_idat;
    end
  end

  function automatic [385:0] MUX_v_386_2_2;
    input [385:0] input_0;
    input [385:0] input_1;
    input  sel;
    reg [385:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_386_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_bbox_req_stream_rsci_bbox_req_stream_wait_ctrl
// ------------------------------------------------------------------


module bbox_core_bbox_req_stream_rsci_bbox_req_stream_wait_ctrl (
  core_wen, bbox_req_stream_rsci_oswt_unreg, bbox_req_stream_rsci_iswt0, bbox_req_stream_rsci_biwt,
      bbox_req_stream_rsci_bdwt, bbox_req_stream_rsci_bcwt, bbox_req_stream_rsci_irdy_core_sct,
      bbox_req_stream_rsci_ivld
);
  input core_wen;
  input bbox_req_stream_rsci_oswt_unreg;
  input bbox_req_stream_rsci_iswt0;
  output bbox_req_stream_rsci_biwt;
  output bbox_req_stream_rsci_bdwt;
  input bbox_req_stream_rsci_bcwt;
  output bbox_req_stream_rsci_irdy_core_sct;
  input bbox_req_stream_rsci_ivld;


  // Interconnect Declarations
  wire bbox_req_stream_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign bbox_req_stream_rsci_bdwt = bbox_req_stream_rsci_oswt_unreg & core_wen;
  assign bbox_req_stream_rsci_biwt = bbox_req_stream_rsci_ogwt & bbox_req_stream_rsci_ivld;
  assign bbox_req_stream_rsci_ogwt = bbox_req_stream_rsci_iswt0 & (~ bbox_req_stream_rsci_bcwt);
  assign bbox_req_stream_rsci_irdy_core_sct = bbox_req_stream_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module ist_core_core_fsm (
  clk, arst_n, core_wen, fsm_output
);
  input clk;
  input arst_n;
  input core_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for ist_core_core_fsm_1
  parameter
    core_rlp_C_0 = 1'd0,
    main_C_0 = 1'd1;

  reg  state_var;
  reg  state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : ist_core_core_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = main_C_0;
      end
      // core_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= core_rlp_C_0;
    end
    else if ( core_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_staller
// ------------------------------------------------------------------


module ist_core_staller (
  clk, arst_n, core_wen, core_wten, ist_req_stream_rsci_wen_comp, ist_resp_stream_rsci_wen_comp,
      core_flen_unreg
);
  input clk;
  input arst_n;
  output core_wen;
  output core_wten;
  input ist_req_stream_rsci_wen_comp;
  input ist_resp_stream_rsci_wen_comp;
  input core_flen_unreg;


  // Interconnect Declarations
  reg core_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign core_wen = ist_req_stream_rsci_wen_comp & ist_resp_stream_rsci_wen_comp
      & (~ core_flen_unreg);
  assign core_wten = core_wten_reg;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      core_wten_reg <= 1'b0;
    end
    else begin
      core_wten_reg <= ~ core_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_28_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_28
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_28_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_28
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_28_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_28_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_28_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_28_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_28_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_28_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_28_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_28_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_28_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_28_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_28_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_28_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_28_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_28_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_28_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_28_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_28_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_28_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_28_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_28_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_28_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_28_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_28_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_28_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_28_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_28_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_28_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_28_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_28_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_28_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_28_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_28_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_28_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_28_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_28_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_28_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_28_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_28
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_28_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_28
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_28_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_28_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_28_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_28_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_28_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_28_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_28_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_28_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_28_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_28_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_28_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_28_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_28_cs_lp_piped_fp_mult_23_8_0_cmp_28_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_28_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_28_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_28_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_28_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_28_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_28_cs_lp_piped_fp_mult_23_8_0_cmp_28_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_28_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_28_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_28_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_28_cs_lp_piped_fp_mult_23_8_0_cmp_28_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_28_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_28_cs_lp_piped_fp_mult_23_8_0_cmp_28_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_28_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_28_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_28_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_28_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_28_cs_lp_piped_fp_mult_23_8_0_cmp_28_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_28_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_1_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_28_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_27_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_27
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_27_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_27
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_27_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_27_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_27_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_27_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_27_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_27_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_27_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_27_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_27_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_27_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_27_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_27_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_27_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_27_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_27_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_27_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_27_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_27_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_27_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_27_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_27_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_27_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_27_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_27_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_27_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_27_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_27_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_27_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_27_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_27_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_27_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_27_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_27_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_27_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_27_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_27_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_27_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_27
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_27_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_27
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_27_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_27_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_27_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_27_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_27_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_27_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_27_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_27_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_27_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_27_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_27_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_27_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_27_cs_lp_piped_fp_mult_23_8_0_cmp_27_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_27_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_27_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_27_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_27_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_27_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_27_cs_lp_piped_fp_mult_23_8_0_cmp_27_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_27_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_27_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_27_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_27_cs_lp_piped_fp_mult_23_8_0_cmp_27_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_27_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_27_cs_lp_piped_fp_mult_23_8_0_cmp_27_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_27_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_27_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_27_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_27_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_27_cs_lp_piped_fp_mult_23_8_0_cmp_27_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_27_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_2_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_27_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_26_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_26
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_26_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_26
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_26_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_26_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_26_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_26_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_26_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_26_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_26_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_26_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_26_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_26_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_26_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_26_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_26_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_26_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_3_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_3_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_26_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_26_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_26_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_26_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_26_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_26_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_26_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_26_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_26_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_26_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_26_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_26_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_26_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_26_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_26_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_26_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_26_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_26_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_3_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_26_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_26_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_3_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_3_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_26_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_3_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_26_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_26_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_26
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_26_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_26
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_26_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_26_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_26_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_26_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_26_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_26_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_26_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_26_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_26_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_26_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_26_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_26_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_26_cs_lp_piped_fp_mult_23_8_0_cmp_26_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_26_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_26_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_3_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_3_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_26_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_26_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_26_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_26_cs_lp_piped_fp_mult_23_8_0_cmp_26_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_26_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_26_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_26_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_26_cs_lp_piped_fp_mult_23_8_0_cmp_26_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_26_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_26_cs_lp_piped_fp_mult_23_8_0_cmp_26_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_26_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_26_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_26_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_3_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_26_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_26_cs_lp_piped_fp_mult_23_8_0_cmp_26_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_3_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_3_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_26_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_3_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_26_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_25_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_25
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_25_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_25
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_25_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_25_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_25_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_25_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_25_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_25_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_25_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_25_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_25_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_25_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_25_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_25_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_25_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_25_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_4_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_4_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_25_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_25_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_25_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_25_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_25_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_25_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_25_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_25_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_25_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_25_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_25_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_25_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_25_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_25_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_25_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_25_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_25_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_25_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_4_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_25_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_25_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_4_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_4_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_25_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_4_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_25_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_25_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_25
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_25_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_25
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_25_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_25_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_25_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_25_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_25_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_25_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_25_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_25_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_25_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_25_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_25_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_25_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_25_cs_lp_piped_fp_mult_23_8_0_cmp_25_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_25_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_25_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_4_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_4_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_25_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_25_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_25_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_25_cs_lp_piped_fp_mult_23_8_0_cmp_25_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_25_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_25_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_25_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_25_cs_lp_piped_fp_mult_23_8_0_cmp_25_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_25_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_25_cs_lp_piped_fp_mult_23_8_0_cmp_25_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_25_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_25_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_25_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_4_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_25_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_25_cs_lp_piped_fp_mult_23_8_0_cmp_25_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_4_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_4_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_25_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_4_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_25_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_24_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_24
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_24_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_24
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_24_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_24_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_24_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_24_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_24_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_24_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_24_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_24_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_24_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_24_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_24_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_24_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_24_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_24_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_5_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_5_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_24_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_24_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_24_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_24_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_24_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_24_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_24_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_24_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_24_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_24_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_24_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_24_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_24_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_24_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_24_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_24_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_24_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_24_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_5_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_24_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_24_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_5_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_5_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_24_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_5_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_24_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_24_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_24
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_24_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_24
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_24_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_24_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_24_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_24_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_24_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_24_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_24_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_24_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_24_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_24_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_24_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_24_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_24_cs_lp_piped_fp_mult_23_8_0_cmp_24_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_24_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_24_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_5_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_5_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_24_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_24_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_24_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_24_cs_lp_piped_fp_mult_23_8_0_cmp_24_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_24_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_24_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_24_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_24_cs_lp_piped_fp_mult_23_8_0_cmp_24_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_24_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_24_cs_lp_piped_fp_mult_23_8_0_cmp_24_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_24_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_24_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_24_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_5_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_24_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_24_cs_lp_piped_fp_mult_23_8_0_cmp_24_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_5_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_5_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_24_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_5_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_24_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_23_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_23
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_23_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_23
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_23_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_23_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_23_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_23_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_23_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_23_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_23_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_23_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_6_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_6_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_23_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_23_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_23_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_23_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_23_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_23_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_23_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_6_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_23_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_23_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_6_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_6_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_23_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_6_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_23_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_23_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_23
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_23_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_23
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_23_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_23_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_23_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_23_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_23_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_23_cs_lp_piped_fp_mult_23_8_0_cmp_23_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_23_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_23_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_6_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_6_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_23_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_23_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_23_cs_lp_piped_fp_mult_23_8_0_cmp_23_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_23_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_23_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_cs_lp_piped_fp_mult_23_8_0_cmp_23_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_cs_lp_piped_fp_mult_23_8_0_cmp_23_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_23_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_6_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_23_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_23_cs_lp_piped_fp_mult_23_8_0_cmp_23_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_6_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_6_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_23_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_6_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_23_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_22
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_22
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_22_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_22_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_22_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_22_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_22_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_22_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_7_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_7_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_22_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_22_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_22_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_22_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_22_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_22_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_22_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_7_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_22_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_22_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_7_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_7_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_22_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_7_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_22_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_22
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_22
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_22_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_22_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_22_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_22_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_22_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_22_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_22_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_22_cs_lp_piped_fp_mult_23_8_0_cmp_22_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_22_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_7_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_7_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_22_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_22_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_22_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_22_cs_lp_piped_fp_mult_23_8_0_cmp_22_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_22_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_22_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_cs_lp_piped_fp_mult_23_8_0_cmp_22_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_cs_lp_piped_fp_mult_23_8_0_cmp_22_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_22_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_7_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_22_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_22_cs_lp_piped_fp_mult_23_8_0_cmp_22_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_7_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_7_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_22_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_7_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_22_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_21_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_21
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_21_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_21
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_21_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_21_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_21_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_21_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_21_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_21_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_21_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_21_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_8_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_8_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_21_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_21_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_21_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_21_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_21_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_21_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_21_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_8_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_21_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_21_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_8_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_8_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_21_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_8_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_21_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_21_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_21
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_21_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_21
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_21_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_21_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_21_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_21_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_21_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_21_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_21_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_21_cs_lp_piped_fp_mult_23_8_0_cmp_21_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_21_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_21_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_8_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_8_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_21_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_21_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_21_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_21_cs_lp_piped_fp_mult_23_8_0_cmp_21_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_21_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_21_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_cs_lp_piped_fp_mult_23_8_0_cmp_21_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_cs_lp_piped_fp_mult_23_8_0_cmp_21_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_21_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_8_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_21_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_21_cs_lp_piped_fp_mult_23_8_0_cmp_21_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_8_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_8_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_21_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_8_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_21_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_20
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_20
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_20_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_20_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_20_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_20_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_20_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_20_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_9_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_9_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_20_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_20_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_20_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_20_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_20_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_20_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_20_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_9_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_20_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_20_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_9_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_9_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_20_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_9_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_20_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_20
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_20
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_20_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_20_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_20_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_20_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_20_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_20_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_20_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_20_cs_lp_piped_fp_mult_23_8_0_cmp_20_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_20_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_9_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_9_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_20_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_20_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_20_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_20_cs_lp_piped_fp_mult_23_8_0_cmp_20_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_20_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_20_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_cs_lp_piped_fp_mult_23_8_0_cmp_20_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_cs_lp_piped_fp_mult_23_8_0_cmp_20_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_20_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_9_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_20_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_20_cs_lp_piped_fp_mult_23_8_0_cmp_20_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_9_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_9_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_20_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_9_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_20_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_19_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_19
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_19_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_19
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_19_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_19_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_19_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_19_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_19_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_19_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_19_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_19_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_10_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_10_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_19_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_19_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_19_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_19_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_19_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_19_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_19_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_10_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_19_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_19_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_10_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_10_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_19_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_10_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_19_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_19_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_19
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_19_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_19
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_19_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_19_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_19_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_19_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_19_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_19_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_19_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_19_cs_lp_piped_fp_mult_23_8_0_cmp_19_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_19_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_19_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_10_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_10_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_19_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_19_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_19_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_19_cs_lp_piped_fp_mult_23_8_0_cmp_19_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_19_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_19_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_cs_lp_piped_fp_mult_23_8_0_cmp_19_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_cs_lp_piped_fp_mult_23_8_0_cmp_19_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_19_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_10_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_19_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_19_cs_lp_piped_fp_mult_23_8_0_cmp_19_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_10_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_10_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_19_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_10_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_19_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_18
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_18
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_18_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_18_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_18_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_18_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_18_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_18_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_11_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_11_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_18_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_18_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_18_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_18_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_18_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_18_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_18_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_11_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_18_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_18_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_11_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_11_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_18_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_11_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_18_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_18
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_18
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_18_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_18_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_18_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_18_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_18_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_18_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_18_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_18_cs_lp_piped_fp_mult_23_8_0_cmp_18_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_18_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_11_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_11_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_18_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_18_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_18_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_18_cs_lp_piped_fp_mult_23_8_0_cmp_18_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_18_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_18_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_cs_lp_piped_fp_mult_23_8_0_cmp_18_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_cs_lp_piped_fp_mult_23_8_0_cmp_18_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_18_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_11_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_18_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_18_cs_lp_piped_fp_mult_23_8_0_cmp_18_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_11_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_11_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_18_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_11_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_18_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_17_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_17
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_17_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_17
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_17_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_17_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_17_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_17_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_17_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_17_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_17_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_17_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_12_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_12_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_17_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_17_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_17_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_17_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_17_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_17_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_17_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_12_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_17_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_17_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_12_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_12_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_17_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_12_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_17_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_17_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_17
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_17_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_17
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_17_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_17_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_17_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_17_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_17_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_17_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_17_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_17_cs_lp_piped_fp_mult_23_8_0_cmp_17_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_17_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_17_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_12_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_12_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_17_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_17_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_17_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_17_cs_lp_piped_fp_mult_23_8_0_cmp_17_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_17_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_17_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_cs_lp_piped_fp_mult_23_8_0_cmp_17_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_cs_lp_piped_fp_mult_23_8_0_cmp_17_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_17_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_12_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_17_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_17_cs_lp_piped_fp_mult_23_8_0_cmp_17_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_12_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_12_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_17_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_12_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_17_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_16
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_16
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_16_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_16_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_16_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_16_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_16_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_16_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_13_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_13_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_16_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_16_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_16_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_16_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_16_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_16_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_16_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_13_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_16_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_16_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_13_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_13_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_16_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_13_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_16_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_16
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_16
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_16_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_16_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_16_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_16_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_16_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_16_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_16_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_16_cs_lp_piped_fp_mult_23_8_0_cmp_16_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_16_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_13_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_13_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_16_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_16_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_16_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_16_cs_lp_piped_fp_mult_23_8_0_cmp_16_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_16_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_16_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_cs_lp_piped_fp_mult_23_8_0_cmp_16_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_cs_lp_piped_fp_mult_23_8_0_cmp_16_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_16_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_13_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_16_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_16_cs_lp_piped_fp_mult_23_8_0_cmp_16_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_13_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_13_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_16_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_13_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_16_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_15_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_15
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_15_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_15
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_15_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_15_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_15_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_15_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_15_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_15_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_15_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_15_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_14_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_14_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_15_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_15_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_15_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_15_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_15_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_15_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_15_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_14_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_15_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_15_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_14_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_14_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_15_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_14_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_15_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_15_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_15
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_15_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_15
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_15_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_15_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_15_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_15_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_15_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_15_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_15_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_15_cs_lp_piped_fp_mult_23_8_0_cmp_15_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_15_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_15_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_14_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_14_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_15_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_15_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_15_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_15_cs_lp_piped_fp_mult_23_8_0_cmp_15_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_15_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_15_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_cs_lp_piped_fp_mult_23_8_0_cmp_15_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_cs_lp_piped_fp_mult_23_8_0_cmp_15_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_15_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_14_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_15_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_15_cs_lp_piped_fp_mult_23_8_0_cmp_15_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_14_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_14_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_15_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_14_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_15_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_14
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_14
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_14_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_14_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_14_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_14_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_14_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_14_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_15_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_15_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_14_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_14_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_14_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_14_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_14_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_14_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_14_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_15_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_14_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_14_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_15_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_15_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_14_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_15_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_14_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_14
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_14
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_14_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_14_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_14_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_14_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_14_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_14_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_14_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_14_cs_lp_piped_fp_mult_23_8_0_cmp_14_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_14_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_15_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_15_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_14_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_14_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_14_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_14_cs_lp_piped_fp_mult_23_8_0_cmp_14_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_14_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_14_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_cs_lp_piped_fp_mult_23_8_0_cmp_14_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_cs_lp_piped_fp_mult_23_8_0_cmp_14_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_14_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_15_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_14_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_14_cs_lp_piped_fp_mult_23_8_0_cmp_14_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_15_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_15_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_14_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_15_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_14_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_13_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_13
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_13_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_13
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_13_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_13_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_13_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_13_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_13_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_13_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_13_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_13_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_16_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_16_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_13_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_13_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_13_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_13_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_13_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_13_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_13_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_16_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_13_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_13_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_16_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_16_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_13_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_16_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_13_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_13_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_13
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_13_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_13
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_13_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_13_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_13_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_13_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_13_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_13_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_13_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_13_cs_lp_piped_fp_mult_23_8_0_cmp_13_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_13_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_13_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_16_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_16_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_13_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_13_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_13_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_13_cs_lp_piped_fp_mult_23_8_0_cmp_13_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_13_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_13_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_cs_lp_piped_fp_mult_23_8_0_cmp_13_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_cs_lp_piped_fp_mult_23_8_0_cmp_13_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_13_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_16_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_13_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_13_cs_lp_piped_fp_mult_23_8_0_cmp_13_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_16_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_16_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_13_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_16_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_13_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_12
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_12
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_12_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_12_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_12_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_12_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_12_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_12_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_17_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_17_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_12_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_12_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_12_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_12_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_12_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_12_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_12_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_17_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_12_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_12_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_17_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_17_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_12_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_17_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_12_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_12
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_12
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_12_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_12_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_12_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_12_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_12_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_12_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_12_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_12_cs_lp_piped_fp_mult_23_8_0_cmp_12_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_12_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_17_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_17_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_12_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_12_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_12_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_12_cs_lp_piped_fp_mult_23_8_0_cmp_12_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_12_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_12_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_cs_lp_piped_fp_mult_23_8_0_cmp_12_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_cs_lp_piped_fp_mult_23_8_0_cmp_12_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_12_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_17_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_12_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_12_cs_lp_piped_fp_mult_23_8_0_cmp_12_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_17_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_17_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_12_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_17_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_12_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_11_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_11
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_11_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_11
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_11_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_11_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_11_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_11_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_11_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_11_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_11_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_11_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_18_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_18_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_11_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_11_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_11_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_11_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_11_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_11_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_11_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_18_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_11_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_11_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_18_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_18_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_11_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_18_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_11_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_11_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_11
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_11_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_11
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_11_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_11_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_11_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_11_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_11_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_11_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_11_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_11_cs_lp_piped_fp_mult_23_8_0_cmp_11_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_11_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_11_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_18_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_18_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_11_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_11_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_11_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_11_cs_lp_piped_fp_mult_23_8_0_cmp_11_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_11_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_11_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_cs_lp_piped_fp_mult_23_8_0_cmp_11_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_cs_lp_piped_fp_mult_23_8_0_cmp_11_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_11_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_18_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_11_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_11_cs_lp_piped_fp_mult_23_8_0_cmp_11_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_18_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_18_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_11_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_18_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_11_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_10
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_10
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_10_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_10_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_10_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_10_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_10_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_10_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_19_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_19_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_10_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_10_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_10_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_10_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_10_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_10_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_10_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_19_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_10_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_10_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_19_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_19_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_10_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_19_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_10_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_10
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_10
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_10_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_10_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_10_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_10_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_10_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_10_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_10_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_10_cs_lp_piped_fp_mult_23_8_0_cmp_10_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_10_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_19_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_19_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_10_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_10_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_10_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_10_cs_lp_piped_fp_mult_23_8_0_cmp_10_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_10_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_10_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_cs_lp_piped_fp_mult_23_8_0_cmp_10_pdswt0
          <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_cs_lp_piped_fp_mult_23_8_0_cmp_10_pdswt0
          <= (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_10_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_19_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_10_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_10_cs_lp_piped_fp_mult_23_8_0_cmp_10_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_19_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_19_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_10_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_19_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_10_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_9_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_9
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_9_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_9
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_9_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_9_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_9_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_9_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_9_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_9_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_9_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_9_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_20_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_20_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_9_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_9_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_9_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_9_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_9_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_9_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_9_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_20_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_9_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_9_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_20_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_20_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_9_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_20_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_9_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_9_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_9
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_9_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_9
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_9_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_9_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_9_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_9_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_9_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_9_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_9_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_9_cs_lp_piped_fp_mult_23_8_0_cmp_9_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_9_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_9_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_20_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_20_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_9_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_9_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_9_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_9_cs_lp_piped_fp_mult_23_8_0_cmp_9_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_9_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_9_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_cs_lp_piped_fp_mult_23_8_0_cmp_9_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_cs_lp_piped_fp_mult_23_8_0_cmp_9_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_9_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_20_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_9_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_9_cs_lp_piped_fp_mult_23_8_0_cmp_9_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_20_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_20_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_9_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_20_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_9_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_8
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_8
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_8_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_8_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_8_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_8_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_8_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_8_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_21_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_21_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_8_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_8_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_8_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_8_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_8_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_8_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_8_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_21_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_8_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_8_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_21_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_21_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_8_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_21_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_8_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_8
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_8
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_8_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_8_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_8_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_8_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_8_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_8_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_8_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_8_cs_lp_piped_fp_mult_23_8_0_cmp_8_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_8_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_21_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_21_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_8_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_8_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_8_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_8_cs_lp_piped_fp_mult_23_8_0_cmp_8_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_8_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_8_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_cs_lp_piped_fp_mult_23_8_0_cmp_8_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_cs_lp_piped_fp_mult_23_8_0_cmp_8_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_8_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_21_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_8_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_8_cs_lp_piped_fp_mult_23_8_0_cmp_8_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_21_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_21_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_8_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_21_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_8_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_7_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_7
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_7_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_7
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_7_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_7_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_7_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_7_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_7_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_7_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_7_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_7_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_22_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_22_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_7_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_7_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_7_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_7_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_7_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_7_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_7_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_22_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_7_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_7_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_22_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_22_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_7_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_22_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_7_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_7_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_7
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_7_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_7
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_7_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_7_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_7_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_7_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_7_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_7_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_7_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_7_cs_lp_piped_fp_mult_23_8_0_cmp_7_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_7_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_7_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_22_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_22_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_7_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_7_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_7_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_7_cs_lp_piped_fp_mult_23_8_0_cmp_7_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_7_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_7_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_cs_lp_piped_fp_mult_23_8_0_cmp_7_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_cs_lp_piped_fp_mult_23_8_0_cmp_7_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_7_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_22_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_7_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_7_cs_lp_piped_fp_mult_23_8_0_cmp_7_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_22_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_22_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_7_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_22_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_7_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_6
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_6
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_6_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_6_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_6_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_6_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_6_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_6_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_23_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_23_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_6_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_6_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_6_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_6_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_6_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_6_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_6_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_23_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_6_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_6_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_23_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_23_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_6_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_23_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_6_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_6
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_6
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_6_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_6_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_6_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_6_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_6_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_6_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_6_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_6_cs_lp_piped_fp_mult_23_8_0_cmp_6_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_6_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_23_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_23_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_6_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_6_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_6_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_6_cs_lp_piped_fp_mult_23_8_0_cmp_6_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_6_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_6_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_cs_lp_piped_fp_mult_23_8_0_cmp_6_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_cs_lp_piped_fp_mult_23_8_0_cmp_6_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_6_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_23_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_6_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_6_cs_lp_piped_fp_mult_23_8_0_cmp_6_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_23_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_23_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_6_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_23_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_6_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_5
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_5
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_5_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_5_a_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_5_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_5_a,
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_5_bawt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_5_a_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_5_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_5_bdwt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_5_a;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_5_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_5_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_5_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_24_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_24_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_5_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_5_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_5_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_5_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_bcwt);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_5_a = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_5_a_core[30:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_5_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_5_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_5_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_24_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_5_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_5_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_24_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_24_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_5_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_24_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_5_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_5
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_5
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_5_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_5_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_5_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_5_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_5_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_5_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_5_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_5_cs_lp_piped_fp_mult_23_8_0_cmp_5_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_5_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_5_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_24_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_24_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_5_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_5_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_5_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_5_cs_lp_piped_fp_mult_23_8_0_cmp_5_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_5_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_5_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_cs_lp_piped_fp_mult_23_8_0_cmp_5_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_cs_lp_piped_fp_mult_23_8_0_cmp_5_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_5_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_24_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_5_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_5_cs_lp_piped_fp_mult_23_8_0_cmp_5_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_24_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_24_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_5_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_24_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_5_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_4
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_4
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_4_a_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_4_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_4_a,
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_a_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_4_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_4_bdwt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_a;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_4_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_25_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_25_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_4_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_4_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_4_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_bcwt);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_4_a = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_4_a_core[30:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_4_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_4_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_4_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_25_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_4_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_4_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_25_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_25_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_4_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_25_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_4_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_4
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_4
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_4_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_4_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_4_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_4_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_4_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_4_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_4_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_4_cs_lp_piped_fp_mult_23_8_0_cmp_4_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_4_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_25_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_25_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_4_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_4_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_4_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_4_cs_lp_piped_fp_mult_23_8_0_cmp_4_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_4_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_4_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_cs_lp_piped_fp_mult_23_8_0_cmp_4_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_cs_lp_piped_fp_mult_23_8_0_cmp_4_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_4_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_25_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_4_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_4_cs_lp_piped_fp_mult_23_8_0_cmp_4_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_25_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_25_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_4_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_25_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_4_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_3_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_3
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_3_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_3
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_3_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_3_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_3_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_3_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_3_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_3_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_3_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_3_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_26_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_26_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_3_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_3_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_3_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_3_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_3_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_3_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_3_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_26_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_3_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_3_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_26_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_26_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_3_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_26_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_3_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_3_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_3
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_3_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_3
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_3_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_3_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_3_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_3_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_3_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_3_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_3_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_3_cs_lp_piped_fp_mult_23_8_0_cmp_3_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_3_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_3_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_26_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_26_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_3_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_3_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_3_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_3_cs_lp_piped_fp_mult_23_8_0_cmp_3_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_3_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_3_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_cs_lp_piped_fp_mult_23_8_0_cmp_3_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_cs_lp_piped_fp_mult_23_8_0_cmp_3_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_3_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_26_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_3_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_3_cs_lp_piped_fp_mult_23_8_0_cmp_3_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_26_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_26_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_3_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_26_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_3_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_2
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_2
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_2_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_27_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_27_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_2_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_2_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_2_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_2_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_27_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_27_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_27_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_2_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_27_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_2_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_2
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_2
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_2_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_2_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_2_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_2_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_2_cs_lp_piped_fp_mult_23_8_0_cmp_2_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_2_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_27_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_27_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_2_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_2_cs_lp_piped_fp_mult_23_8_0_cmp_2_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_2_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_2_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_cs_lp_piped_fp_mult_23_8_0_cmp_2_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_cs_lp_piped_fp_mult_23_8_0_cmp_2_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_2_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_27_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_2_cs_lp_piped_fp_mult_23_8_0_cmp_2_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_27_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_27_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_2_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_27_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_2_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_1
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_1
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_1_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_28_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_28_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_1_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_1_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_1_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_1_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_28_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_28_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_28_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_1_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_28_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_1_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_1
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_1
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_1_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt, ccs_lp_piped_fp_mult_23_8_0_cmp_1_launch_core_sct,
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_1_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_1_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_1_cs_lp_piped_fp_mult_23_8_0_cmp_1_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_1_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_28_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_28_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_1_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_1_cs_lp_piped_fp_mult_23_8_0_cmp_1_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_1_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_1_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_cs_lp_piped_fp_mult_23_8_0_cmp_1_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_cs_lp_piped_fp_mult_23_8_0_cmp_1_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_1_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_28_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_1_cs_lp_piped_fp_mult_23_8_0_cmp_1_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_28_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_28_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_1_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_28_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_1_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp
    (
  clk, arst_n, ccs_lp_piped_fp_mult_23_8_0_cmp_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_bawt;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_biwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_bcwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_z_bfwt_1;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_bawt = ccs_lp_piped_fp_mult_23_8_0_cmp_biwt
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_bcwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_mult_23_8_0_cmp_z,
      ccs_lp_piped_fp_mult_23_8_0_cmp_z_bfwt, ccs_lp_piped_fp_mult_23_8_0_cmp_z_bfwt_1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_bcwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_mult_23_8_0_cmp_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_mult_23_8_0_cmp_biwt ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_z_bfwt <= ccs_lp_piped_fp_mult_23_8_0_cmp_z;
      ccs_lp_piped_fp_mult_23_8_0_cmp_z_bfwt_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_biwt);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_1_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_bcwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_1_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_oswt_unreg, ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_biwt, ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_launch_core_sct, ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_oswt_unreg;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_biwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_launch_core_sct;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_cs_lp_piped_fp_mult_23_8_0_cmp_pdswt0;
  reg [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_mult_23_8_0_cmp_icwt;

  wire[1:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_nl;
  wire[2:0] nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt = ccs_lp_piped_fp_mult_23_8_0_cmp_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_biwt = ccs_lp_piped_fp_mult_23_8_0_cmp_cs_lp_piped_fp_mult_23_8_0_cmp_pdswt0
      | (ccs_lp_piped_fp_mult_23_8_0_cmp_icwt!=2'b00);
  assign ccs_lp_piped_fp_mult_23_8_0_cmp_launch_core_sct = core_wen & ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_cs_lp_piped_fp_mult_23_8_0_cmp_pdswt0 <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_mult_23_8_0_cmp_cs_lp_piped_fp_mult_23_8_0_cmp_pdswt0 <= (~
          core_wten) & ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1;
      ccs_lp_piped_fp_mult_23_8_0_cmp_icwt <= nl_ccs_lp_piped_fp_mult_23_8_0_cmp_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_mult_23_8_0_cmp_cs_lp_piped_fp_mult_23_8_0_cmp_pdswt0);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_nl = nl_lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_mult_23_8_0_cmp_icwt  = lp_piped_fp_mult_AC_RND_CONV_0_32_8_acc_nl
      + ccs_lp_piped_fp_mult_23_8_0_cmp_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_17_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_17
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_17_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_17
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_17_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_17_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_17_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_17_bdwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_17_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_17_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_17_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_17_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_17_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_17_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_17_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_17_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_17_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_17_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_17_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_17_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_17_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_17_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_17_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_17_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_17_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_17_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_17_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_17_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_17_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_17_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_17_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_17_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_17_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_17_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_17_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_17_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_17_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_17_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_17_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_17_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_17_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_17
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_17_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_17
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_17_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_17_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_17_biwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_17_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_17_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_17_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_17_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_17_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_17_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_17_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_17_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_17_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_17_cs_lp_piped_fp_add_23_8_0_cmp_17_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_17_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_17_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_17_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_17_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_17_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_17_cs_lp_piped_fp_add_23_8_0_cmp_17_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_17_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_17_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_17_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_17_cs_lp_piped_fp_add_23_8_0_cmp_17_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_17_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_17_cs_lp_piped_fp_add_23_8_0_cmp_17_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_add_23_8_0_cmp_17_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_17_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_17_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_17_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_17_cs_lp_piped_fp_add_23_8_0_cmp_17_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_17_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_1_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_17_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_16_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_16
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_16_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_16
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_16_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_16_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_16_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_16_bdwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_16_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_16_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_16_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_16_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_16_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_16_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_16_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_16_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_16_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_16_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_16_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_16_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_16_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_16_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_16_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_16_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_16_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_16_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_16_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_16_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_16_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_16_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_16_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_16_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_16_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_16_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_16_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_16_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_16_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_16_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_16_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_16_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_16_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_16
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_16_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_16
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_16_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_16_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_16_biwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_16_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_16_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_16_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_16_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_16_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_16_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_16_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_16_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_16_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_16_cs_lp_piped_fp_add_23_8_0_cmp_16_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_16_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_16_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_16_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_16_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_16_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_16_cs_lp_piped_fp_add_23_8_0_cmp_16_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_16_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_16_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_16_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_16_cs_lp_piped_fp_add_23_8_0_cmp_16_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_16_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_16_cs_lp_piped_fp_add_23_8_0_cmp_16_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_add_23_8_0_cmp_16_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_16_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_16_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_16_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_16_cs_lp_piped_fp_add_23_8_0_cmp_16_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_16_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_2_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_16_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_15_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_15
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_15_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_15
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_15_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_15_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_15_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_15_bdwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_15_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_15_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_15_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_15_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_15_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_15_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_15_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_15_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_15_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_15_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_3_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_3_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_15_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_15_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_15_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_15_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_15_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_15_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_15_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_15_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_15_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_15_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_15_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_15_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_15_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_15_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_15_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_15_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_15_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_15_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_3_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_15_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_15_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_3_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_3_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_15_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_3_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_15_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_15_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_15
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_15_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_15
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_15_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_15_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_15_biwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_15_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_15_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_15_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_15_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_15_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_15_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_15_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_15_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_15_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_15_cs_lp_piped_fp_add_23_8_0_cmp_15_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_15_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_15_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_3_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_3_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_15_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_15_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_15_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_15_cs_lp_piped_fp_add_23_8_0_cmp_15_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_15_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_15_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_15_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_15_cs_lp_piped_fp_add_23_8_0_cmp_15_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_15_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_15_cs_lp_piped_fp_add_23_8_0_cmp_15_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_add_23_8_0_cmp_15_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_15_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_15_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_3_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_15_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_15_cs_lp_piped_fp_add_23_8_0_cmp_15_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_3_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_3_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_15_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_3_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_15_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_14_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_14
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_14_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_14
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_14_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_14_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_14_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_14_bdwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_14_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_14_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_14_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_14_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_14_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_14_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_14_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_14_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_14_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_14_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_4_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_4_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_14_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_14_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_14_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_14_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_14_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_14_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_14_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_14_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_14_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_14_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_14_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_14_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_14_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_14_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_14_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_14_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_14_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_14_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_4_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_14_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_14_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_4_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_4_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_14_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_4_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_14_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_14_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_14
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_14_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_14
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_14_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_14_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_14_biwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_14_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_14_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_14_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_14_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_14_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_14_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_14_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_14_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_14_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_14_cs_lp_piped_fp_add_23_8_0_cmp_14_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_14_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_14_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_4_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_4_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_14_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_14_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_14_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_14_cs_lp_piped_fp_add_23_8_0_cmp_14_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_14_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_14_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_14_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_14_cs_lp_piped_fp_add_23_8_0_cmp_14_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_14_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_14_cs_lp_piped_fp_add_23_8_0_cmp_14_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_add_23_8_0_cmp_14_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_14_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_14_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_4_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_14_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_14_cs_lp_piped_fp_add_23_8_0_cmp_14_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_4_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_4_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_14_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_4_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_14_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_13_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_13
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_13_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_13
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_13_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_13_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_13_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_13_bdwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_13_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_13_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_13_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_13_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_13_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_13_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_13_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_13_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_13_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_13_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_5_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_5_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_13_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_13_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_13_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_13_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_13_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_13_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_13_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_13_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_13_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_13_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_13_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_13_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_13_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_13_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_13_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_13_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_13_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_13_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_5_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_13_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_13_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_5_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_5_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_13_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_5_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_13_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_13_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_13
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_13_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_13
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_13_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_13_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_13_biwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_13_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_13_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_13_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_13_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_13_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_13_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_13_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_13_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_13_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_13_cs_lp_piped_fp_add_23_8_0_cmp_13_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_13_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_13_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_5_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_5_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_13_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_13_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_13_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_13_cs_lp_piped_fp_add_23_8_0_cmp_13_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_13_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_13_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_13_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_13_cs_lp_piped_fp_add_23_8_0_cmp_13_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_13_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_13_cs_lp_piped_fp_add_23_8_0_cmp_13_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_add_23_8_0_cmp_13_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_13_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_13_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_5_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_13_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_13_cs_lp_piped_fp_add_23_8_0_cmp_13_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_5_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_5_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_13_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_5_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_13_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_12_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_12
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_12_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_12
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_12_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_12_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_12_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_12_bdwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_12_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_12_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_12_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_12_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_12_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_12_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_12_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_12_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_12_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_12_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_6_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_6_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_12_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_12_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_12_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_12_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_12_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_12_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_12_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_12_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_12_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_12_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_12_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_12_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_12_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_12_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_12_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_12_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_12_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_12_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_6_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_12_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_12_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_6_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_6_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_12_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_6_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_12_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_12_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_12
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_12_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_12
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_12_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_12_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_12_biwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_12_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_12_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_12_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_12_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_12_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_12_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_12_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_12_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_12_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_12_cs_lp_piped_fp_add_23_8_0_cmp_12_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_12_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_12_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_6_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_6_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_12_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_12_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_12_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_12_cs_lp_piped_fp_add_23_8_0_cmp_12_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_12_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_12_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_12_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_12_cs_lp_piped_fp_add_23_8_0_cmp_12_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_12_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_12_cs_lp_piped_fp_add_23_8_0_cmp_12_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_add_23_8_0_cmp_12_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_12_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_12_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_6_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_12_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_12_cs_lp_piped_fp_add_23_8_0_cmp_12_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_6_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_6_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_12_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_6_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_12_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_11_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_11
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_11_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_11
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_11_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_11_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_11_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_11_bdwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_11_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_11_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_11_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_11_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_11_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_11_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_11_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_11_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_11_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_11_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_7_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_7_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_11_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_11_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_11_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_11_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_11_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_11_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_11_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_11_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_11_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_11_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_11_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_11_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_11_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_11_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_11_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_11_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_11_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_11_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_7_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_11_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_11_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_7_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_7_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_11_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_7_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_11_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_11_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_11
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_11_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_11
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_11_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_11_biwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_11_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_11_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_11_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_11_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_11_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_11_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_11_cs_lp_piped_fp_add_23_8_0_cmp_11_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_11_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_11_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_7_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_7_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_11_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_11_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_11_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_11_cs_lp_piped_fp_add_23_8_0_cmp_11_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_11_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_11_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_11_cs_lp_piped_fp_add_23_8_0_cmp_11_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_11_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_11_cs_lp_piped_fp_add_23_8_0_cmp_11_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_11_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_11_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_7_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_11_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_11_cs_lp_piped_fp_add_23_8_0_cmp_11_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_7_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_7_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_11_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_7_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_11_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_10_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_10
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_10_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_10
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_10_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_10_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_10_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_10_bdwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_10_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_10_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_10_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_10_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_10_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_10_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_10_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_10_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_10_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_10_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_8_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_8_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_10_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_10_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_10_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_10_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_10_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_10_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_10_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_10_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_10_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_10_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_10_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_10_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_10_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_10_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_10_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_10_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_10_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_10_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_8_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_10_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_10_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_8_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_8_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_10_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_8_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_10_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_10_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_10
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_10_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_10
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_10_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_10_biwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_10_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_10_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_10_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_10_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_10_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_10_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_10_cs_lp_piped_fp_add_23_8_0_cmp_10_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_10_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_10_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_8_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_8_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_10_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_10_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_10_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_10_cs_lp_piped_fp_add_23_8_0_cmp_10_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_10_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_10_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_10_cs_lp_piped_fp_add_23_8_0_cmp_10_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_10_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_10_cs_lp_piped_fp_add_23_8_0_cmp_10_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_10_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_10_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_8_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_10_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_10_cs_lp_piped_fp_add_23_8_0_cmp_10_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_8_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_8_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_10_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_8_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_10_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_9_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_9
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_9_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_9
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_9_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_9_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_9_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_9_bdwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_9_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_9_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_9_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_9_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_9_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_9_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_9_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_9_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_9_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_9_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_9_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_9_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_9_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_9_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_9_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_9_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_9_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_9_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_9_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_9_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_9_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_9_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_9_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_9_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_9_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_9_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_9_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_9_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_9_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_9_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_9_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_9_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_9_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_9_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_9_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_9_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_9_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_9_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_9_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_9
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_9_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_9
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_9_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_9_biwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_9_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_9_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_9_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_9_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_9_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_9_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_9_cs_lp_piped_fp_add_23_8_0_cmp_9_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_9_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_9_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_9_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_9_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_9_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_9_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_9_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_9_cs_lp_piped_fp_add_23_8_0_cmp_9_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_9_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_9_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_9_cs_lp_piped_fp_add_23_8_0_cmp_9_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_9_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_9_cs_lp_piped_fp_add_23_8_0_cmp_9_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_9_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_9_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_9_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_9_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_9_cs_lp_piped_fp_add_23_8_0_cmp_9_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_9_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_9_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_9_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_9_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_9_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_8_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_8
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_8_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_8
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_8_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_8_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_8_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_8_bdwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_8_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_8_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_8_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_8_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_8_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_8_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_8_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_8_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_8_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_8_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_10_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_10_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_8_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_8_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_8_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_8_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_8_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_8_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_8_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_8_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_8_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_8_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_8_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_8_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_8_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_8_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_8_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_8_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_8_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_8_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_10_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_8_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_8_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_10_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_10_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_8_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_10_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_8_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_8_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_8
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_8_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_8
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_8_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_8_biwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_8_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_8_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_8_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_8_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_8_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_8_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_8_cs_lp_piped_fp_add_23_8_0_cmp_8_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_8_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_8_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_10_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_10_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_8_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_8_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_8_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_8_cs_lp_piped_fp_add_23_8_0_cmp_8_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_8_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_8_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_8_cs_lp_piped_fp_add_23_8_0_cmp_8_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_8_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_8_cs_lp_piped_fp_add_23_8_0_cmp_8_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_8_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_8_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_10_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_8_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_8_cs_lp_piped_fp_add_23_8_0_cmp_8_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_10_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_10_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_8_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_10_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_8_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_7_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_7
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_7_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_7
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_7_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_7_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_7_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_7_bdwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_7_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_7_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_7_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_7_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_7_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_7_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_7_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_7_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_7_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_7_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_11_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_11_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_7_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_7_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_7_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_7_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_7_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_7_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_7_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_7_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_7_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_7_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_7_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_7_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_7_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_7_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_7_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_7_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_7_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_7_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_11_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_7_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_7_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_11_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_11_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_7_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_11_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_7_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_7_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_7
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_7_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_7
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_7_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_7_biwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_7_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_7_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_7_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_7_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_7_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_7_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_7_cs_lp_piped_fp_add_23_8_0_cmp_7_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_7_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_7_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_11_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_11_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_7_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_7_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_7_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_7_cs_lp_piped_fp_add_23_8_0_cmp_7_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_7_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_7_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_7_cs_lp_piped_fp_add_23_8_0_cmp_7_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_7_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_7_cs_lp_piped_fp_add_23_8_0_cmp_7_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_7_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_7_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_11_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_7_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_7_cs_lp_piped_fp_add_23_8_0_cmp_7_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_11_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_11_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_7_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_11_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_7_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_6_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_6
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_6_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_6
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_6_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_6_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_6_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_6_bdwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_6_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_6_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_6_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_6_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_6_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_6_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_6_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_6_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_6_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_6_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_12_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_12_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_6_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_6_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_6_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_6_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_6_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_6_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_6_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_6_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_6_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_6_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_6_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_6_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_6_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_6_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_6_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_6_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_6_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_6_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_12_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_6_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_6_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_12_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_12_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_6_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_12_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_6_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_6_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_6
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_6_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_6
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_6_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_6_biwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_6_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_6_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_6_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_6_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_6_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_6_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_6_cs_lp_piped_fp_add_23_8_0_cmp_6_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_6_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_6_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_12_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_12_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_6_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_6_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_6_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_6_cs_lp_piped_fp_add_23_8_0_cmp_6_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_6_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_6_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_6_cs_lp_piped_fp_add_23_8_0_cmp_6_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_6_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_6_cs_lp_piped_fp_add_23_8_0_cmp_6_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_6_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_6_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_12_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_6_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_6_cs_lp_piped_fp_add_23_8_0_cmp_6_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_12_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_12_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_6_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_12_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_6_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_5_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_5
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_5_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_5
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_5_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_5_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_5_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_5_bdwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_5_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_5_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_5_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_5_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_5_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_5_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_5_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_5_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_5_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_5_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_13_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_13_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_5_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_5_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_5_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_5_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_5_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_5_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_5_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_5_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_5_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_5_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_5_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_5_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_5_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_5_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_5_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_5_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_5_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_5_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_13_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_5_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_5_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_13_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_13_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_5_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_13_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_5_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_5_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_5
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_5_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_5
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_5_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_5_biwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_5_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_5_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_5_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_5_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_5_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_5_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_5_cs_lp_piped_fp_add_23_8_0_cmp_5_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_5_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_5_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_13_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_13_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_5_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_5_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_5_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_5_cs_lp_piped_fp_add_23_8_0_cmp_5_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_5_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_5_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_5_cs_lp_piped_fp_add_23_8_0_cmp_5_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_5_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_5_cs_lp_piped_fp_add_23_8_0_cmp_5_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_5_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_5_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_13_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_5_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_5_cs_lp_piped_fp_add_23_8_0_cmp_5_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_13_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_13_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_5_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_13_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_5_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_4_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_4
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_4_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_4
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_4_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_4_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_4_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_4_bdwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_4_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_4_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_4_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_4_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_4_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_4_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_4_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_4_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_4_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_4_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_14_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_14_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_4_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_4_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_4_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_4_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_4_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_4_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_4_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_4_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_4_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_4_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_4_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_4_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_4_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_4_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_4_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_4_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_4_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_4_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_14_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_4_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_4_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_14_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_14_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_4_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_14_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_4_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_4_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_4
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_4_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_4
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_4_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_4_biwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_4_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_4_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_4_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_4_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_4_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_4_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_4_cs_lp_piped_fp_add_23_8_0_cmp_4_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_4_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_4_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_14_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_14_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_4_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_4_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_4_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_4_cs_lp_piped_fp_add_23_8_0_cmp_4_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_4_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_4_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_4_cs_lp_piped_fp_add_23_8_0_cmp_4_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_4_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_4_cs_lp_piped_fp_add_23_8_0_cmp_4_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_4_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_4_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_14_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_4_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_4_cs_lp_piped_fp_add_23_8_0_cmp_4_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_14_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_14_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_4_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_14_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_4_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_3_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_3
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_3_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_3
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_3_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_3_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_3_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_3_bdwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_3_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_3_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_3_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_3_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_3_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_3_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_3_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_3_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_3_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_3_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_15_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_15_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_3_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_3_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_3_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_3_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_3_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_3_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_3_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_3_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_3_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_3_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_3_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_3_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_3_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_3_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_3_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_3_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_3_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_3_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_15_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_3_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_3_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_15_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_15_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_3_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_15_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_3_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_3_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_3
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_3_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_3
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_3_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_3_biwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_3_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_3_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_3_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_3_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_3_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_3_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_3_cs_lp_piped_fp_add_23_8_0_cmp_3_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_3_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_3_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_15_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_15_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_3_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_3_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_3_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_3_cs_lp_piped_fp_add_23_8_0_cmp_3_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_3_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_3_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_3_cs_lp_piped_fp_add_23_8_0_cmp_3_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_3_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_3_cs_lp_piped_fp_add_23_8_0_cmp_3_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_3_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_3_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_15_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_3_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_3_cs_lp_piped_fp_add_23_8_0_cmp_3_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_15_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_15_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_3_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_15_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_3_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_2
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_2
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_2_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_2_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_16_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_16_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_2_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_2_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_2_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_2_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_2_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_2_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_2_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_2_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_2_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_2_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_2_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_2_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_2_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_2_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_16_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_16_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_16_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_2_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_16_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_2_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_2
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_2
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_2_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_2_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_2_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_2_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_2_cs_lp_piped_fp_add_23_8_0_cmp_2_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_2_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_16_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_16_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_2_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_2_cs_lp_piped_fp_add_23_8_0_cmp_2_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_2_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_2_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_2_cs_lp_piped_fp_add_23_8_0_cmp_2_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_2_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_2_cs_lp_piped_fp_add_23_8_0_cmp_2_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_2_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_2_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_16_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_2_cs_lp_piped_fp_add_23_8_0_cmp_2_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_16_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_16_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_2_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_16_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_2_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_1
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_1
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_1_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_1_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_17_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_17_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_1_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_1_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_1_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_1_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_1_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_1_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_1_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_1_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_1_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_1_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_1_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_1_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_1_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_1_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_17_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_17_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_17_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_1_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_17_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_1_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_1
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_1
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_1_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_1_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_1_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_1_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_1_cs_lp_piped_fp_add_23_8_0_cmp_1_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_1_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_17_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_17_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_1_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_1_cs_lp_piped_fp_add_23_8_0_cmp_1_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_1_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_1_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_1_cs_lp_piped_fp_add_23_8_0_cmp_1_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_1_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_1_cs_lp_piped_fp_add_23_8_0_cmp_1_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_1_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_1_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_17_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_1_cs_lp_piped_fp_add_23_8_0_cmp_1_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_17_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_17_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_1_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_17_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_1_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp
    (
  clk, arst_n, ccs_lp_piped_fp_add_23_8_0_cmp_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_add_23_8_0_cmp_bawt;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_biwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_bdwt;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_bcwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_z_bfwt_1;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_bawt = ccs_lp_piped_fp_add_23_8_0_cmp_biwt
      | (ccs_lp_piped_fp_add_23_8_0_cmp_bcwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_add_23_8_0_cmp_z,
      ccs_lp_piped_fp_add_23_8_0_cmp_z_bfwt, ccs_lp_piped_fp_add_23_8_0_cmp_z_bfwt_1,
      ccs_lp_piped_fp_add_23_8_0_cmp_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_bcwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_add_23_8_0_cmp_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_add_23_8_0_cmp_biwt ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_z_bfwt <= ccs_lp_piped_fp_add_23_8_0_cmp_z;
      ccs_lp_piped_fp_add_23_8_0_cmp_z_bfwt_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_biwt);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_1_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_bcwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_1_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_oswt_unreg, ccs_lp_piped_fp_add_23_8_0_cmp_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_biwt, ccs_lp_piped_fp_add_23_8_0_cmp_bdwt, ccs_lp_piped_fp_add_23_8_0_cmp_launch_core_sct,
      ccs_lp_piped_fp_add_23_8_0_cmp_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_oswt_unreg;
  input ccs_lp_piped_fp_add_23_8_0_cmp_iswt1;
  output ccs_lp_piped_fp_add_23_8_0_cmp_biwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_bdwt;
  output ccs_lp_piped_fp_add_23_8_0_cmp_launch_core_sct;
  input ccs_lp_piped_fp_add_23_8_0_cmp_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_add_23_8_0_cmp_cs_lp_piped_fp_add_23_8_0_cmp_pdswt0;
  reg [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_add_23_8_0_cmp_icwt;

  wire[1:0] lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_nl;
  wire[2:0] nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_add_23_8_0_cmp_bdwt = ccs_lp_piped_fp_add_23_8_0_cmp_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_add_23_8_0_cmp_biwt = ccs_lp_piped_fp_add_23_8_0_cmp_cs_lp_piped_fp_add_23_8_0_cmp_pdswt0
      | (ccs_lp_piped_fp_add_23_8_0_cmp_icwt!=2'b00);
  assign ccs_lp_piped_fp_add_23_8_0_cmp_launch_core_sct = core_wen & ccs_lp_piped_fp_add_23_8_0_cmp_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_cs_lp_piped_fp_add_23_8_0_cmp_pdswt0 <= 1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_add_23_8_0_cmp_cs_lp_piped_fp_add_23_8_0_cmp_pdswt0 <= (~ core_wten)
          & ccs_lp_piped_fp_add_23_8_0_cmp_iswt1;
      ccs_lp_piped_fp_add_23_8_0_cmp_icwt <= nl_ccs_lp_piped_fp_add_23_8_0_cmp_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_add_23_8_0_cmp_cs_lp_piped_fp_add_23_8_0_cmp_pdswt0);
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_nl = nl_lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_add_23_8_0_cmp_icwt  = lp_piped_fp_add_AC_RND_CONV_0_32_8_acc_nl
      + ccs_lp_piped_fp_add_23_8_0_cmp_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_recip_23_8_0_cmp_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_dp
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_recip_23_8_0_cmp_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_dp
    (
  clk, arst_n, ccs_lp_piped_fp_recip_23_8_0_cmp_bawt, ccs_lp_piped_fp_recip_23_8_0_cmp_a_core,
      ccs_lp_piped_fp_recip_23_8_0_cmp_z_mxwt, ccs_lp_piped_fp_recip_23_8_0_cmp_biwt,
      ccs_lp_piped_fp_recip_23_8_0_cmp_bdwt, ccs_lp_piped_fp_recip_23_8_0_cmp_a,
      ccs_lp_piped_fp_recip_23_8_0_cmp_z
);
  input clk;
  input arst_n;
  output ccs_lp_piped_fp_recip_23_8_0_cmp_bawt;
  input [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_a_core;
  output [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_z_mxwt;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_biwt;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_bdwt;
  output [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_a;
  input [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_z;


  // Interconnect Declarations
  reg [1:0] ccs_lp_piped_fp_recip_23_8_0_cmp_bcwt;
  wire [2:0] nl_ccs_lp_piped_fp_recip_23_8_0_cmp_bcwt;
  reg [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_z_bfwt;
  reg [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_z_bfwt_1;

  wire[1:0] lp_piped_fp_recip_AC_RND_CONV_0_32_8_acc_1_nl;
  wire[2:0] nl_lp_piped_fp_recip_AC_RND_CONV_0_32_8_acc_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_recip_23_8_0_cmp_bawt = ccs_lp_piped_fp_recip_23_8_0_cmp_biwt
      | (ccs_lp_piped_fp_recip_23_8_0_cmp_bcwt!=2'b00);
  assign ccs_lp_piped_fp_recip_23_8_0_cmp_z_mxwt = MUX_v_32_3_2(ccs_lp_piped_fp_recip_23_8_0_cmp_z,
      ccs_lp_piped_fp_recip_23_8_0_cmp_z_bfwt, ccs_lp_piped_fp_recip_23_8_0_cmp_z_bfwt_1,
      ccs_lp_piped_fp_recip_23_8_0_cmp_bcwt);
  assign ccs_lp_piped_fp_recip_23_8_0_cmp_a = {1'b0 , (ccs_lp_piped_fp_recip_23_8_0_cmp_a_core[30:0])};
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_recip_23_8_0_cmp_bcwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_recip_23_8_0_cmp_bcwt <= nl_ccs_lp_piped_fp_recip_23_8_0_cmp_bcwt[1:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_recip_23_8_0_cmp_z_bfwt <= 32'b00000000000000000000000000000000;
      ccs_lp_piped_fp_recip_23_8_0_cmp_z_bfwt_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( ccs_lp_piped_fp_recip_23_8_0_cmp_biwt ) begin
      ccs_lp_piped_fp_recip_23_8_0_cmp_z_bfwt <= ccs_lp_piped_fp_recip_23_8_0_cmp_z;
      ccs_lp_piped_fp_recip_23_8_0_cmp_z_bfwt_1 <= ccs_lp_piped_fp_recip_23_8_0_cmp_z_bfwt;
    end
  end
  assign nl_lp_piped_fp_recip_AC_RND_CONV_0_32_8_acc_1_nl = conv_s2s_1_2(ccs_lp_piped_fp_recip_23_8_0_cmp_bdwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_recip_23_8_0_cmp_biwt);
  assign lp_piped_fp_recip_AC_RND_CONV_0_32_8_acc_1_nl = nl_lp_piped_fp_recip_AC_RND_CONV_0_32_8_acc_1_nl[1:0];
  assign nl_ccs_lp_piped_fp_recip_23_8_0_cmp_bcwt  = lp_piped_fp_recip_AC_RND_CONV_0_32_8_acc_1_nl
      + ccs_lp_piped_fp_recip_23_8_0_cmp_bcwt;

  function automatic [31:0] MUX_v_32_3_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [31:0] input_2;
    input [1:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = input_0;
      end
      2'b01 : begin
        result = input_1;
      end
      default : begin
        result = input_2;
      end
    endcase
    MUX_v_32_3_2 = result;
  end
  endfunction


  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_recip_23_8_0_cmp_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_ctrl
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_recip_23_8_0_cmp_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_ctrl
    (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_recip_23_8_0_cmp_oswt_unreg,
      ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1, ccs_lp_piped_fp_recip_23_8_0_cmp_biwt,
      ccs_lp_piped_fp_recip_23_8_0_cmp_bdwt, ccs_lp_piped_fp_recip_23_8_0_cmp_launch_core_sct,
      ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_oswt_unreg;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1;
  output ccs_lp_piped_fp_recip_23_8_0_cmp_biwt;
  output ccs_lp_piped_fp_recip_23_8_0_cmp_bdwt;
  output ccs_lp_piped_fp_recip_23_8_0_cmp_launch_core_sct;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1_pff;


  // Interconnect Declarations
  reg ccs_lp_piped_fp_recip_23_8_0_cmp_cs_lp_piped_fp_recip_23_8_0_cmp_pdswt0;
  reg [1:0] ccs_lp_piped_fp_recip_23_8_0_cmp_icwt;
  wire [2:0] nl_ccs_lp_piped_fp_recip_23_8_0_cmp_icwt;

  wire[1:0] lp_piped_fp_recip_AC_RND_CONV_0_32_8_acc_nl;
  wire[2:0] nl_lp_piped_fp_recip_AC_RND_CONV_0_32_8_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ccs_lp_piped_fp_recip_23_8_0_cmp_bdwt = ccs_lp_piped_fp_recip_23_8_0_cmp_oswt_unreg
      & core_wen;
  assign ccs_lp_piped_fp_recip_23_8_0_cmp_biwt = ccs_lp_piped_fp_recip_23_8_0_cmp_cs_lp_piped_fp_recip_23_8_0_cmp_pdswt0
      | (ccs_lp_piped_fp_recip_23_8_0_cmp_icwt!=2'b00);
  assign ccs_lp_piped_fp_recip_23_8_0_cmp_launch_core_sct = core_wen & ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1_pff;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_recip_23_8_0_cmp_cs_lp_piped_fp_recip_23_8_0_cmp_pdswt0 <=
          1'b0;
      ccs_lp_piped_fp_recip_23_8_0_cmp_icwt <= 2'b00;
    end
    else begin
      ccs_lp_piped_fp_recip_23_8_0_cmp_cs_lp_piped_fp_recip_23_8_0_cmp_pdswt0 <=
          (~ core_wten) & ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1;
      ccs_lp_piped_fp_recip_23_8_0_cmp_icwt <= nl_ccs_lp_piped_fp_recip_23_8_0_cmp_icwt[1:0];
    end
  end
  assign nl_lp_piped_fp_recip_AC_RND_CONV_0_32_8_acc_nl = conv_s2s_1_2(ccs_lp_piped_fp_recip_23_8_0_cmp_biwt)
      + conv_u2s_1_2(ccs_lp_piped_fp_recip_23_8_0_cmp_cs_lp_piped_fp_recip_23_8_0_cmp_pdswt0);
  assign lp_piped_fp_recip_AC_RND_CONV_0_32_8_acc_nl = nl_lp_piped_fp_recip_AC_RND_CONV_0_32_8_acc_nl[1:0];
  assign nl_ccs_lp_piped_fp_recip_23_8_0_cmp_icwt  = lp_piped_fp_recip_AC_RND_CONV_0_32_8_acc_nl
      + ccs_lp_piped_fp_recip_23_8_0_cmp_icwt;

  function automatic [1:0] conv_s2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_s2s_1_2 = {vector[0], vector};
  end
  endfunction


  function automatic [1:0] conv_u2s_1_2 ;
    input [0:0]  vector ;
  begin
    conv_u2s_1_2 =  {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ist_resp_stream_rsci_ist_resp_stream_wait_dp
// ------------------------------------------------------------------


module ist_core_ist_resp_stream_rsci_ist_resp_stream_wait_dp (
  clk, arst_n, ist_resp_stream_rsci_oswt_unreg, ist_resp_stream_rsci_bawt, ist_resp_stream_rsci_wen_comp,
      ist_resp_stream_rsci_biwt, ist_resp_stream_rsci_bdwt, ist_resp_stream_rsci_bcwt
);
  input clk;
  input arst_n;
  input ist_resp_stream_rsci_oswt_unreg;
  output ist_resp_stream_rsci_bawt;
  output ist_resp_stream_rsci_wen_comp;
  input ist_resp_stream_rsci_biwt;
  input ist_resp_stream_rsci_bdwt;
  output ist_resp_stream_rsci_bcwt;
  reg ist_resp_stream_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign ist_resp_stream_rsci_bawt = ist_resp_stream_rsci_biwt | ist_resp_stream_rsci_bcwt;
  assign ist_resp_stream_rsci_wen_comp = (~ ist_resp_stream_rsci_oswt_unreg) | ist_resp_stream_rsci_bawt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ist_resp_stream_rsci_bcwt <= 1'b0;
    end
    else begin
      ist_resp_stream_rsci_bcwt <= ~((~(ist_resp_stream_rsci_bcwt | ist_resp_stream_rsci_biwt))
          | ist_resp_stream_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ist_resp_stream_rsci_ist_resp_stream_wait_ctrl
// ------------------------------------------------------------------


module ist_core_ist_resp_stream_rsci_ist_resp_stream_wait_ctrl (
  core_wen, ist_resp_stream_rsci_oswt_unreg, ist_resp_stream_rsci_iswt0, ist_resp_stream_rsci_biwt,
      ist_resp_stream_rsci_bdwt, ist_resp_stream_rsci_bcwt, ist_resp_stream_rsci_irdy,
      ist_resp_stream_rsci_ivld_core_sct
);
  input core_wen;
  input ist_resp_stream_rsci_oswt_unreg;
  input ist_resp_stream_rsci_iswt0;
  output ist_resp_stream_rsci_biwt;
  output ist_resp_stream_rsci_bdwt;
  input ist_resp_stream_rsci_bcwt;
  input ist_resp_stream_rsci_irdy;
  output ist_resp_stream_rsci_ivld_core_sct;


  // Interconnect Declarations
  wire ist_resp_stream_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign ist_resp_stream_rsci_bdwt = ist_resp_stream_rsci_oswt_unreg & core_wen;
  assign ist_resp_stream_rsci_biwt = ist_resp_stream_rsci_ogwt & ist_resp_stream_rsci_irdy;
  assign ist_resp_stream_rsci_ogwt = ist_resp_stream_rsci_iswt0 & (~ ist_resp_stream_rsci_bcwt);
  assign ist_resp_stream_rsci_ivld_core_sct = ist_resp_stream_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ist_req_stream_rsci_ist_req_stream_wait_dp
// ------------------------------------------------------------------


module ist_core_ist_req_stream_rsci_ist_req_stream_wait_dp (
  clk, arst_n, ist_req_stream_rsci_oswt_unreg, ist_req_stream_rsci_bawt, ist_req_stream_rsci_wen_comp,
      ist_req_stream_rsci_idat_mxwt, ist_req_stream_rsci_biwt, ist_req_stream_rsci_bdwt,
      ist_req_stream_rsci_bcwt, ist_req_stream_rsci_idat
);
  input clk;
  input arst_n;
  input ist_req_stream_rsci_oswt_unreg;
  output ist_req_stream_rsci_bawt;
  output ist_req_stream_rsci_wen_comp;
  output [553:0] ist_req_stream_rsci_idat_mxwt;
  input ist_req_stream_rsci_biwt;
  input ist_req_stream_rsci_bdwt;
  output ist_req_stream_rsci_bcwt;
  reg ist_req_stream_rsci_bcwt;
  input [553:0] ist_req_stream_rsci_idat;


  // Interconnect Declarations
  reg [553:0] ist_req_stream_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign ist_req_stream_rsci_bawt = ist_req_stream_rsci_biwt | ist_req_stream_rsci_bcwt;
  assign ist_req_stream_rsci_wen_comp = (~ ist_req_stream_rsci_oswt_unreg) | ist_req_stream_rsci_bawt;
  assign ist_req_stream_rsci_idat_mxwt = MUX_v_554_2_2(ist_req_stream_rsci_idat,
      ist_req_stream_rsci_idat_bfwt, ist_req_stream_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ist_req_stream_rsci_bcwt <= 1'b0;
    end
    else begin
      ist_req_stream_rsci_bcwt <= ~((~(ist_req_stream_rsci_bcwt | ist_req_stream_rsci_biwt))
          | ist_req_stream_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ist_req_stream_rsci_idat_bfwt <= 554'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ist_req_stream_rsci_biwt ) begin
      ist_req_stream_rsci_idat_bfwt <= ist_req_stream_rsci_idat;
    end
  end

  function automatic [553:0] MUX_v_554_2_2;
    input [553:0] input_0;
    input [553:0] input_1;
    input  sel;
    reg [553:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_554_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ist_req_stream_rsci_ist_req_stream_wait_ctrl
// ------------------------------------------------------------------


module ist_core_ist_req_stream_rsci_ist_req_stream_wait_ctrl (
  core_wen, ist_req_stream_rsci_oswt_unreg, ist_req_stream_rsci_iswt0, ist_req_stream_rsci_biwt,
      ist_req_stream_rsci_bdwt, ist_req_stream_rsci_bcwt, ist_req_stream_rsci_irdy_core_sct,
      ist_req_stream_rsci_ivld
);
  input core_wen;
  input ist_req_stream_rsci_oswt_unreg;
  input ist_req_stream_rsci_iswt0;
  output ist_req_stream_rsci_biwt;
  output ist_req_stream_rsci_bdwt;
  input ist_req_stream_rsci_bcwt;
  output ist_req_stream_rsci_irdy_core_sct;
  input ist_req_stream_rsci_ivld;


  // Interconnect Declarations
  wire ist_req_stream_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign ist_req_stream_rsci_bdwt = ist_req_stream_rsci_oswt_unreg & core_wen;
  assign ist_req_stream_rsci_biwt = ist_req_stream_rsci_ogwt & ist_req_stream_rsci_ivld;
  assign ist_req_stream_rsci_ogwt = ist_req_stream_rsci_iswt0 & (~ ist_req_stream_rsci_bcwt);
  assign ist_req_stream_rsci_irdy_core_sct = ist_req_stream_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_2
// ------------------------------------------------------------------


module init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_2 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_recip_23_8_0_cmp_2_oswt_unreg,
      ccs_lp_piped_fp_recip_23_8_0_cmp_2_bawt, ccs_lp_piped_fp_recip_23_8_0_cmp_2_iswt1,
      ccs_lp_piped_fp_recip_23_8_0_cmp_2_a_core, ccs_lp_piped_fp_recip_23_8_0_cmp_2_z_mxwt,
      ccs_lp_piped_fp_recip_23_8_0_cmp_2_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_2_oswt_unreg;
  output ccs_lp_piped_fp_recip_23_8_0_cmp_2_bawt;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_2_iswt1;
  input [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_2_a_core;
  output [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_2_z_mxwt;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_2_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_2_biwt;
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_2_bdwt;
  wire [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_2_z;
  wire [7:0] ccs_lp_piped_fp_recip_23_8_0_cmp_2_status;
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_2_launch_core_sct;
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_2_pipe_full;
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_2_pipe_ovf;
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_2_arrive;
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_2_push_out_n;
  wire [1:0] ccs_lp_piped_fp_recip_23_8_0_cmp_2_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_recip_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_recip_23_8_0_cmp_2 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_recip_23_8_0_cmp_2_a_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_recip_23_8_0_cmp_2_z),
      .status(ccs_lp_piped_fp_recip_23_8_0_cmp_2_status),
      .launch(ccs_lp_piped_fp_recip_23_8_0_cmp_2_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_recip_23_8_0_cmp_2_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_recip_23_8_0_cmp_2_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_recip_23_8_0_cmp_2_arrive),
      .push_out_n(ccs_lp_piped_fp_recip_23_8_0_cmp_2_push_out_n),
      .pipe_census(ccs_lp_piped_fp_recip_23_8_0_cmp_2_pipe_census)
    );
  init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_2_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_ctrl_2
      init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_2_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_ctrl_2_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_2_oswt_unreg(ccs_lp_piped_fp_recip_23_8_0_cmp_2_oswt_unreg),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_2_iswt1(ccs_lp_piped_fp_recip_23_8_0_cmp_2_iswt1),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_2_biwt(ccs_lp_piped_fp_recip_23_8_0_cmp_2_biwt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_2_bdwt(ccs_lp_piped_fp_recip_23_8_0_cmp_2_bdwt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_2_launch_core_sct(ccs_lp_piped_fp_recip_23_8_0_cmp_2_launch_core_sct),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_2_iswt1_pff(ccs_lp_piped_fp_recip_23_8_0_cmp_2_iswt1_pff)
    );
  init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_2_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_dp_2
      init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_2_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_dp_2_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_2_bawt(ccs_lp_piped_fp_recip_23_8_0_cmp_2_bawt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_2_z_mxwt(ccs_lp_piped_fp_recip_23_8_0_cmp_2_z_mxwt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_2_biwt(ccs_lp_piped_fp_recip_23_8_0_cmp_2_biwt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_2_bdwt(ccs_lp_piped_fp_recip_23_8_0_cmp_2_bdwt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_2_z(ccs_lp_piped_fp_recip_23_8_0_cmp_2_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_1
// ------------------------------------------------------------------


module init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_1 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_recip_23_8_0_cmp_1_oswt_unreg,
      ccs_lp_piped_fp_recip_23_8_0_cmp_1_bawt, ccs_lp_piped_fp_recip_23_8_0_cmp_1_iswt1,
      ccs_lp_piped_fp_recip_23_8_0_cmp_1_a_core, ccs_lp_piped_fp_recip_23_8_0_cmp_1_z_mxwt,
      ccs_lp_piped_fp_recip_23_8_0_cmp_1_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_1_oswt_unreg;
  output ccs_lp_piped_fp_recip_23_8_0_cmp_1_bawt;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_1_iswt1;
  input [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_1_a_core;
  output [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_1_z_mxwt;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_1_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_1_biwt;
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_1_bdwt;
  wire [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_1_z;
  wire [7:0] ccs_lp_piped_fp_recip_23_8_0_cmp_1_status;
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_1_launch_core_sct;
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_1_pipe_full;
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_1_pipe_ovf;
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_1_arrive;
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_1_push_out_n;
  wire [1:0] ccs_lp_piped_fp_recip_23_8_0_cmp_1_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_recip_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_recip_23_8_0_cmp_1 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_recip_23_8_0_cmp_1_a_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_recip_23_8_0_cmp_1_z),
      .status(ccs_lp_piped_fp_recip_23_8_0_cmp_1_status),
      .launch(ccs_lp_piped_fp_recip_23_8_0_cmp_1_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_recip_23_8_0_cmp_1_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_recip_23_8_0_cmp_1_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_recip_23_8_0_cmp_1_arrive),
      .push_out_n(ccs_lp_piped_fp_recip_23_8_0_cmp_1_push_out_n),
      .pipe_census(ccs_lp_piped_fp_recip_23_8_0_cmp_1_pipe_census)
    );
  init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_1_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_ctrl_1
      init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_1_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_ctrl_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_1_oswt_unreg(ccs_lp_piped_fp_recip_23_8_0_cmp_1_oswt_unreg),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_1_iswt1(ccs_lp_piped_fp_recip_23_8_0_cmp_1_iswt1),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_1_biwt(ccs_lp_piped_fp_recip_23_8_0_cmp_1_biwt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_1_bdwt(ccs_lp_piped_fp_recip_23_8_0_cmp_1_bdwt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_1_launch_core_sct(ccs_lp_piped_fp_recip_23_8_0_cmp_1_launch_core_sct),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_1_iswt1_pff(ccs_lp_piped_fp_recip_23_8_0_cmp_1_iswt1_pff)
    );
  init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_1_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_dp_1
      init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_1_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_dp_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_1_bawt(ccs_lp_piped_fp_recip_23_8_0_cmp_1_bawt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_1_z_mxwt(ccs_lp_piped_fp_recip_23_8_0_cmp_1_z_mxwt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_1_biwt(ccs_lp_piped_fp_recip_23_8_0_cmp_1_biwt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_1_bdwt(ccs_lp_piped_fp_recip_23_8_0_cmp_1_bdwt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_1_z(ccs_lp_piped_fp_recip_23_8_0_cmp_1_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_ccs_lp_piped_fp_recip_23_8_0_cmp
// ------------------------------------------------------------------


module init_core_ccs_lp_piped_fp_recip_23_8_0_cmp (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_recip_23_8_0_cmp_oswt_unreg,
      ccs_lp_piped_fp_recip_23_8_0_cmp_bawt, ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1,
      ccs_lp_piped_fp_recip_23_8_0_cmp_a_core, ccs_lp_piped_fp_recip_23_8_0_cmp_z_mxwt,
      ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_oswt_unreg;
  output ccs_lp_piped_fp_recip_23_8_0_cmp_bawt;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1;
  input [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_a_core;
  output [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_z_mxwt;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_biwt;
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_bdwt;
  wire [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_z;
  wire [7:0] ccs_lp_piped_fp_recip_23_8_0_cmp_status;
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_launch_core_sct;
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_pipe_full;
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_pipe_ovf;
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_arrive;
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_push_out_n;
  wire [1:0] ccs_lp_piped_fp_recip_23_8_0_cmp_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_recip_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_recip_23_8_0_cmp (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_recip_23_8_0_cmp_a_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_recip_23_8_0_cmp_z),
      .status(ccs_lp_piped_fp_recip_23_8_0_cmp_status),
      .launch(ccs_lp_piped_fp_recip_23_8_0_cmp_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_recip_23_8_0_cmp_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_recip_23_8_0_cmp_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_recip_23_8_0_cmp_arrive),
      .push_out_n(ccs_lp_piped_fp_recip_23_8_0_cmp_push_out_n),
      .pipe_census(ccs_lp_piped_fp_recip_23_8_0_cmp_pipe_census)
    );
  init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_ctrl
      init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_ctrl_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_oswt_unreg(ccs_lp_piped_fp_recip_23_8_0_cmp_oswt_unreg),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1(ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_biwt(ccs_lp_piped_fp_recip_23_8_0_cmp_biwt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_bdwt(ccs_lp_piped_fp_recip_23_8_0_cmp_bdwt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_launch_core_sct(ccs_lp_piped_fp_recip_23_8_0_cmp_launch_core_sct),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1_pff(ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1_pff)
    );
  init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_dp
      init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_bawt(ccs_lp_piped_fp_recip_23_8_0_cmp_bawt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_z_mxwt(ccs_lp_piped_fp_recip_23_8_0_cmp_z_mxwt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_biwt(ccs_lp_piped_fp_recip_23_8_0_cmp_biwt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_bdwt(ccs_lp_piped_fp_recip_23_8_0_cmp_bdwt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_z(ccs_lp_piped_fp_recip_23_8_0_cmp_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_ccs_lp_piped_fp_add_23_8_0_cmp_2
// ------------------------------------------------------------------


module init_core_ccs_lp_piped_fp_add_23_8_0_cmp_2 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_2_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_2_a_core, ccs_lp_piped_fp_add_23_8_0_cmp_2_b_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt, ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_2_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_2_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_2_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_2_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_2_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_2_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp_2 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_2_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_2_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_2_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_2_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_2_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_2_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_2_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_2_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_2_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_2_pipe_census)
    );
  init_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_2
      init_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_2_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_2_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_2_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1_pff)
    );
  init_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_2
      init_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_2_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_z(ccs_lp_piped_fp_add_23_8_0_cmp_2_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_ccs_lp_piped_fp_add_23_8_0_cmp_1
// ------------------------------------------------------------------


module init_core_ccs_lp_piped_fp_add_23_8_0_cmp_1 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_1_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_1_a_core, ccs_lp_piped_fp_add_23_8_0_cmp_1_b_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt, ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_1_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_1_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_1_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_1_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_1_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_1_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp_1 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_1_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_1_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_1_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_1_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_1_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_1_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_1_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_1_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_1_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_1_pipe_census)
    );
  init_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_1
      init_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_1_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_1_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1_pff)
    );
  init_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_1
      init_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_z(ccs_lp_piped_fp_add_23_8_0_cmp_1_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_ccs_lp_piped_fp_add_23_8_0_cmp
// ------------------------------------------------------------------


module init_core_ccs_lp_piped_fp_add_23_8_0_cmp (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_oswt_unreg, ccs_lp_piped_fp_add_23_8_0_cmp_bawt,
      ccs_lp_piped_fp_add_23_8_0_cmp_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_a_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_b_core, ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_pipe_census)
    );
  init_core_ccs_lp_piped_fp_add_23_8_0_cmp_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl
      init_core_ccs_lp_piped_fp_add_23_8_0_cmp_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_iswt1_pff)
    );
  init_core_ccs_lp_piped_fp_add_23_8_0_cmp_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp
      init_core_ccs_lp_piped_fp_add_23_8_0_cmp_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_z(ccs_lp_piped_fp_add_23_8_0_cmp_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2
// ------------------------------------------------------------------


module init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_2_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_2_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_2_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_2_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_2_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_2_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_2_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_2_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_2 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_2_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_2_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_2_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_2_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_2_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_2_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_2_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_2_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_2_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_2_pipe_census)
    );
  init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_2
      init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_2_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_2_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_2_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1_pff)
    );
  init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_2
      init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_2_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_z(ccs_lp_piped_fp_mult_23_8_0_cmp_2_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1
// ------------------------------------------------------------------


module init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_1_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_1_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_1_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_1_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_1_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_1_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_1_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_1_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_1 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_1_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_1_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_1_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_1_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_1_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_1_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_1_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_1_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_1_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_1_pipe_census)
    );
  init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_1
      init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_1_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_1_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1_pff)
    );
  init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_1
      init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_z(ccs_lp_piped_fp_mult_23_8_0_cmp_1_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_ccs_lp_piped_fp_mult_23_8_0_cmp
// ------------------------------------------------------------------


module init_core_ccs_lp_piped_fp_mult_23_8_0_cmp (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_oswt_unreg, ccs_lp_piped_fp_mult_23_8_0_cmp_bawt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_a_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_b_core, ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_pipe_census)
    );
  init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl
      init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1_pff)
    );
  init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp
      init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_z(ccs_lp_piped_fp_mult_23_8_0_cmp_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_trv_req_stream_rsci
// ------------------------------------------------------------------


module init_core_trv_req_stream_rsci (
  clk, arst_n, trv_req_stream_rsc_dat, trv_req_stream_rsc_vld, trv_req_stream_rsc_rdy,
      core_wen, trv_req_stream_rsci_oswt_unreg, trv_req_stream_rsci_bawt, trv_req_stream_rsci_iswt0,
      trv_req_stream_rsci_wen_comp, trv_req_stream_rsci_idat
);
  input clk;
  input arst_n;
  output [457:0] trv_req_stream_rsc_dat;
  output trv_req_stream_rsc_vld;
  input trv_req_stream_rsc_rdy;
  input core_wen;
  input trv_req_stream_rsci_oswt_unreg;
  output trv_req_stream_rsci_bawt;
  input trv_req_stream_rsci_iswt0;
  output trv_req_stream_rsci_wen_comp;
  input [457:0] trv_req_stream_rsci_idat;


  // Interconnect Declarations
  wire trv_req_stream_rsci_biwt;
  wire trv_req_stream_rsci_bdwt;
  wire trv_req_stream_rsci_bcwt;
  wire trv_req_stream_rsci_irdy;
  wire trv_req_stream_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd17),
  .width(32'sd458)) trv_req_stream_rsci (
      .irdy(trv_req_stream_rsci_irdy),
      .ivld(trv_req_stream_rsci_ivld_core_sct),
      .idat(trv_req_stream_rsci_idat),
      .rdy(trv_req_stream_rsc_rdy),
      .vld(trv_req_stream_rsc_vld),
      .dat(trv_req_stream_rsc_dat)
    );
  init_core_trv_req_stream_rsci_trv_req_stream_wait_ctrl init_core_trv_req_stream_rsci_trv_req_stream_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .trv_req_stream_rsci_oswt_unreg(trv_req_stream_rsci_oswt_unreg),
      .trv_req_stream_rsci_iswt0(trv_req_stream_rsci_iswt0),
      .trv_req_stream_rsci_biwt(trv_req_stream_rsci_biwt),
      .trv_req_stream_rsci_bdwt(trv_req_stream_rsci_bdwt),
      .trv_req_stream_rsci_bcwt(trv_req_stream_rsci_bcwt),
      .trv_req_stream_rsci_irdy(trv_req_stream_rsci_irdy),
      .trv_req_stream_rsci_ivld_core_sct(trv_req_stream_rsci_ivld_core_sct)
    );
  init_core_trv_req_stream_rsci_trv_req_stream_wait_dp init_core_trv_req_stream_rsci_trv_req_stream_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .trv_req_stream_rsci_oswt_unreg(trv_req_stream_rsci_oswt_unreg),
      .trv_req_stream_rsci_bawt(trv_req_stream_rsci_bawt),
      .trv_req_stream_rsci_wen_comp(trv_req_stream_rsci_wen_comp),
      .trv_req_stream_rsci_biwt(trv_req_stream_rsci_biwt),
      .trv_req_stream_rsci_bdwt(trv_req_stream_rsci_bdwt),
      .trv_req_stream_rsci_bcwt(trv_req_stream_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core_init_req_stream_rsci
// ------------------------------------------------------------------


module init_core_init_req_stream_rsci (
  clk, arst_n, init_req_stream_rsc_dat, init_req_stream_rsc_vld, init_req_stream_rsc_rdy,
      core_wen, init_req_stream_rsci_oswt_unreg, init_req_stream_rsci_bawt, init_req_stream_rsci_iswt0,
      init_req_stream_rsci_wen_comp, init_req_stream_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [361:0] init_req_stream_rsc_dat;
  input init_req_stream_rsc_vld;
  output init_req_stream_rsc_rdy;
  input core_wen;
  input init_req_stream_rsci_oswt_unreg;
  output init_req_stream_rsci_bawt;
  input init_req_stream_rsci_iswt0;
  output init_req_stream_rsci_wen_comp;
  output [361:0] init_req_stream_rsci_idat_mxwt;


  // Interconnect Declarations
  wire init_req_stream_rsci_biwt;
  wire init_req_stream_rsci_bdwt;
  wire init_req_stream_rsci_bcwt;
  wire init_req_stream_rsci_irdy_core_sct;
  wire init_req_stream_rsci_ivld;
  wire [361:0] init_req_stream_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd16),
  .width(32'sd362)) init_req_stream_rsci (
      .rdy(init_req_stream_rsc_rdy),
      .vld(init_req_stream_rsc_vld),
      .dat(init_req_stream_rsc_dat),
      .irdy(init_req_stream_rsci_irdy_core_sct),
      .ivld(init_req_stream_rsci_ivld),
      .idat(init_req_stream_rsci_idat)
    );
  init_core_init_req_stream_rsci_init_req_stream_wait_ctrl init_core_init_req_stream_rsci_init_req_stream_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .init_req_stream_rsci_oswt_unreg(init_req_stream_rsci_oswt_unreg),
      .init_req_stream_rsci_iswt0(init_req_stream_rsci_iswt0),
      .init_req_stream_rsci_biwt(init_req_stream_rsci_biwt),
      .init_req_stream_rsci_bdwt(init_req_stream_rsci_bdwt),
      .init_req_stream_rsci_bcwt(init_req_stream_rsci_bcwt),
      .init_req_stream_rsci_irdy_core_sct(init_req_stream_rsci_irdy_core_sct),
      .init_req_stream_rsci_ivld(init_req_stream_rsci_ivld)
    );
  init_core_init_req_stream_rsci_init_req_stream_wait_dp init_core_init_req_stream_rsci_init_req_stream_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .init_req_stream_rsci_oswt_unreg(init_req_stream_rsci_oswt_unreg),
      .init_req_stream_rsci_bawt(init_req_stream_rsci_bawt),
      .init_req_stream_rsci_wen_comp(init_req_stream_rsci_wen_comp),
      .init_req_stream_rsci_idat_mxwt(init_req_stream_rsci_idat_mxwt),
      .init_req_stream_rsci_biwt(init_req_stream_rsci_biwt),
      .init_req_stream_rsci_bdwt(init_req_stream_rsci_bdwt),
      .init_req_stream_rsci_bcwt(init_req_stream_rsci_bcwt),
      .init_req_stream_rsci_idat(init_req_stream_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_23
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_23 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_23_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_23_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_23_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_23_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_23_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_23_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_23_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_23_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_23_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_23_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_23_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_23_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_23_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_23_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_23 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_23_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_23_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_23_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_23_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_23_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_23_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_23_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_23_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_23_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_23_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_23_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_23
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_23_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_23_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_23_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_23_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_23_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_23_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_23
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_23_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_23_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_23_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_23_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_23_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_z(ccs_lp_piped_fp_mult_23_8_0_cmp_23_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_22_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_22_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_22_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_22_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_22_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_22_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_a;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_b;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_22_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_22_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_22_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_22_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_22_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_22_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_22_a_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_22_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_22_a_core
      = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_22_a_core[30:16]) , 16'b0000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_22_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_22_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_22_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_22_b_core
      = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_22_b_core[30:23]) , 23'b00000000000000000000000};
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_22 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_22_a),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_22_b),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_22_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_22_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_22_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_22_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_22_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_22_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_22_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_22_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_22
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_22_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_22_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_22_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_22_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_22_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_22
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_22_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_22_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_22_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_22_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_b_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_22_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_22_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_22_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_22_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_a(ccs_lp_piped_fp_mult_23_8_0_cmp_22_a),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_b(ccs_lp_piped_fp_mult_23_8_0_cmp_22_b),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_z(ccs_lp_piped_fp_mult_23_8_0_cmp_22_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_21
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_21 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_21_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_21_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_21_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_21_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_21_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_21_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_21_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_21_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_21_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_21_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_21_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_21_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_21_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_21_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_21_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_21_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_21 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_21_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_21_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_21_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_21_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_21_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_21_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_21_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_21_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_21_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_21_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_21_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_21
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_21_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_21_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_21_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_21_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_21_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_21_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_21_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_21
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_21_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_21_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_21_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_21_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_21_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_z(ccs_lp_piped_fp_mult_23_8_0_cmp_21_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_20_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_20_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_20_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_20_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_20_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_20_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_a;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_b;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_20_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_20_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_20_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_20_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_20_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_20_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_20_a_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_20_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_20_a_core
      = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_20_a_core[30:16]) , 16'b0000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_20_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_20_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_20_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_20_b_core
      = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_20_b_core[30:23]) , 23'b00000000000000000000000};
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_20 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_20_a),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_20_b),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_20_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_20_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_20_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_20_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_20_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_20_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_20_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_20_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_20
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_20_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_20_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_20_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_20_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_20_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_20
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_20_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_20_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_20_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_20_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_b_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_20_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_20_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_20_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_20_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_a(ccs_lp_piped_fp_mult_23_8_0_cmp_20_a),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_b(ccs_lp_piped_fp_mult_23_8_0_cmp_20_b),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_z(ccs_lp_piped_fp_mult_23_8_0_cmp_20_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_19
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_19 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_19_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_19_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_19_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_19_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_19_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_19_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_19_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_19_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_19_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_19_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_19_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_19_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_19_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_19_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_19_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_19_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_19 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_19_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_19_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_19_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_19_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_19_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_19_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_19_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_19_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_19_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_19_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_19_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_19
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_19_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_19_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_19_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_19_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_19_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_19_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_19_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_19
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_19_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_19_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_19_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_19_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_19_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_z(ccs_lp_piped_fp_mult_23_8_0_cmp_19_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_18_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_18_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_18_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_18_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_18_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_18_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_a;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_b;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_18_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_18_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_18_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_18_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_18_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_18_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_18_a_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_18_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_18_a_core
      = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_18_a_core[30:16]) , 16'b0000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_18_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_18_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_18_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_18_b_core
      = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_18_b_core[30:23]) , 23'b00000000000000000000000};
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_18 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_18_a),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_18_b),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_18_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_18_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_18_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_18_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_18_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_18_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_18_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_18_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_18
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_18_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_18_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_18_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_18_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_18_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_18
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_18_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_18_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_18_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_18_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_b_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_18_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_18_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_18_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_18_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_a(ccs_lp_piped_fp_mult_23_8_0_cmp_18_a),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_b(ccs_lp_piped_fp_mult_23_8_0_cmp_18_b),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_z(ccs_lp_piped_fp_mult_23_8_0_cmp_18_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_17
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_17 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_17_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_17_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_17_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_17_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_17_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_17_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_17_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_17_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_17_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_17_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_17_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_17_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_17_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_17_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_17_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_17_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_17 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_17_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_17_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_17_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_17_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_17_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_17_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_17_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_17_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_17_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_17_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_17_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_17
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_17_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_17_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_17_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_17_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_17_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_17_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_17_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_17
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_17_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_17_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_17_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_17_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_17_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_z(ccs_lp_piped_fp_mult_23_8_0_cmp_17_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_16_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_16_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_16_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_16_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_16_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_16_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_a;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_b;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_16_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_16_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_16_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_16_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_16_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_16_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_16_a_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_16_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_16_a_core
      = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_16_a_core[30:16]) , 16'b0000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_16_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_16_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_16_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_16_b_core
      = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_16_b_core[30:23]) , 23'b00000000000000000000000};
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_16 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_16_a),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_16_b),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_16_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_16_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_16_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_16_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_16_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_16_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_16_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_16_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_16
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_16_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_16_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_16_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_16_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_16_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_16
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_16_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_16_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_16_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_16_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_b_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_16_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_16_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_16_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_16_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_a(ccs_lp_piped_fp_mult_23_8_0_cmp_16_a),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_b(ccs_lp_piped_fp_mult_23_8_0_cmp_16_b),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_z(ccs_lp_piped_fp_mult_23_8_0_cmp_16_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_15
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_15 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_15_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_15_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_15_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_15_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_15_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_15_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_15_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_15_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_15_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_15_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_15_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_15_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_15_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_15_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_15_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_15_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_15 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_15_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_15_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_15_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_15_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_15_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_15_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_15_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_15_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_15_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_15_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_15_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_15
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_15_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_15_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_15_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_15_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_15_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_15_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_15_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_15
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_15_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_15_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_15_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_15_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_15_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_z(ccs_lp_piped_fp_mult_23_8_0_cmp_15_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_14_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_14_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_14_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_14_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_14_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_14_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_a;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_b;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_14_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_14_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_14_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_14_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_14_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_14_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_14_a_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_14_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_14_a_core
      = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_14_a_core[30:16]) , 16'b0000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_14_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_14_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_14_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_14_b_core
      = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_14_b_core[30:23]) , 23'b00000000000000000000000};
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_14 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_14_a),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_14_b),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_14_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_14_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_14_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_14_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_14_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_14_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_14_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_14_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_14
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_14_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_14_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_14_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_14_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_14_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_14
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_14_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_14_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_14_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_14_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_b_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_14_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_14_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_14_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_14_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_a(ccs_lp_piped_fp_mult_23_8_0_cmp_14_a),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_b(ccs_lp_piped_fp_mult_23_8_0_cmp_14_b),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_z(ccs_lp_piped_fp_mult_23_8_0_cmp_14_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_13
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_13 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_13_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_13_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_13_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_13_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_13_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_13_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_13_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_13_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_13_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_13_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_13_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_13_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_13_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_13_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_13_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_13_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_13 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_13_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_13_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_13_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_13_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_13_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_13_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_13_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_13_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_13_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_13_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_13_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_13
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_13_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_13_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_13_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_13_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_13_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_13_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_13_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_13
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_13_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_13_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_13_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_13_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_13_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_z(ccs_lp_piped_fp_mult_23_8_0_cmp_13_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_12_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_12_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_12_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_12_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_12_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_12_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_a;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_b;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_12_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_12_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_12_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_12_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_12_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_12_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_12_a_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_12_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_12_a_core
      = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_12_a_core[30:16]) , 16'b0000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_12_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_12_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_12_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_12_b_core
      = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_12_b_core[30:23]) , 23'b00000000000000000000000};
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_12 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_12_a),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_12_b),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_12_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_12_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_12_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_12_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_12_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_12_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_12_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_12_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_12
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_12_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_12_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_12_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_12_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_12_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_12
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_12_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_12_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_12_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_12_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_b_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_12_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_12_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_12_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_12_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_a(ccs_lp_piped_fp_mult_23_8_0_cmp_12_a),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_b(ccs_lp_piped_fp_mult_23_8_0_cmp_12_b),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_z(ccs_lp_piped_fp_mult_23_8_0_cmp_12_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_11
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_11 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_11_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_11_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_11_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_11_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_11_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_11_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_11_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_11_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_11_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_11_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_11_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_11_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_11_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_11_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_11_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_11_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_11 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_11_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_11_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_11_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_11_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_11_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_11_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_11_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_11_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_11_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_11_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_11_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_11
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_11_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_11_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_11_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_11_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_11_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_11_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_11_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_11
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_11_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_11_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_11_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_11_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_11_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_z(ccs_lp_piped_fp_mult_23_8_0_cmp_11_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_10_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_10_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_10_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_10_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_10_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_10_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_a;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_b;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_10_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_10_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_10_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_10_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_10_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_10_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_10_a_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_10_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_10_a_core
      = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_10_a_core[30:16]) , 16'b0000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_10_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_10_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_10_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_10_b_core
      = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_10_b_core[30:23]) , 23'b00000000000000000000000};
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_10 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_10_a),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_10_b),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_10_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_10_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_10_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_10_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_10_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_10_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_10_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_10_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_10
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_10_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_10_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_10_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_10_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_10_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_10
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_10_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_10_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_10_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_10_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_b_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_10_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_10_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_10_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_10_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_a(ccs_lp_piped_fp_mult_23_8_0_cmp_10_a),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_b(ccs_lp_piped_fp_mult_23_8_0_cmp_10_b),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_z(ccs_lp_piped_fp_mult_23_8_0_cmp_10_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_9
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_9 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_9_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_9_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_9_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_9_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_9_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_9_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_9_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_9_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_9_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_9_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_9_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_9_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_9_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_9_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_9_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_9_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_9 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_9_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_9_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_9_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_9_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_9_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_9_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_9_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_9_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_9_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_9_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_9_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_9
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_9_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_9_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_9_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_9_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_9_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_9_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_9_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_9
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_9_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_9_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_9_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_9_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_9_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_z(ccs_lp_piped_fp_mult_23_8_0_cmp_9_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_8_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_8_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_8_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_8_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_8_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_8_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_a;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_b;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_8_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_8_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_8_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_8_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_8_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_8_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_8_a_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_8_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_8_a_core
      = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_8_a_core[30:16]) , 16'b0000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_8_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_8_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_8_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_8_b_core
      = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_8_b_core[30:23]) , 23'b00000000000000000000000};
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_8 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_8_a),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_8_b),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_8_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_8_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_8_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_8_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_8_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_8_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_8_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_8_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_8
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_8_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_8_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_8_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_8_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_8_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_8
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_8_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_8_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_8_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_8_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_b_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_8_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_8_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_8_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_8_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_a(ccs_lp_piped_fp_mult_23_8_0_cmp_8_a),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_b(ccs_lp_piped_fp_mult_23_8_0_cmp_8_b),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_z(ccs_lp_piped_fp_mult_23_8_0_cmp_8_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_7
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_7 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_7_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_7_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_7_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_7_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_7_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_7_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_7_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_7_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_7_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_7_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_7_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_7_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_7_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_7_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_7_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_7_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_7 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_7_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_7_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_7_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_7_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_7_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_7_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_7_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_7_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_7_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_7_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_7_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_7
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_7_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_7_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_7_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_7_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_7_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_7_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_7_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_7
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_7_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_7_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_7_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_7_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_7_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_z(ccs_lp_piped_fp_mult_23_8_0_cmp_7_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_6_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_6_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_6_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_6_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_6_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_6_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_a;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_b;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_6_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_6_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_6_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_6_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_6_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_6_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_6_a_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_6_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_6_a_core
      = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_6_a_core[30:16]) , 16'b0000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_6_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_6_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_6_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_6_b_core
      = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_6_b_core[30:23]) , 23'b00000000000000000000000};
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_6 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_6_a),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_6_b),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_6_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_6_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_6_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_6_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_6_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_6_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_6_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_6_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_6
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_6_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_6_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_6_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_6_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_6_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_6
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_6_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_6_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_6_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_6_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_b_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_6_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_6_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_6_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_6_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_a(ccs_lp_piped_fp_mult_23_8_0_cmp_6_a),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_b(ccs_lp_piped_fp_mult_23_8_0_cmp_6_b),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_z(ccs_lp_piped_fp_mult_23_8_0_cmp_6_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_5_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_5_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_5_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_5_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_5_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_5_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_5_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_5_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_5_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_5_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_5_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_5_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_5_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_5_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_5_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_5_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_5 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_5_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_5_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_5_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_5_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_5_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_5_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_5_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_5_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_5_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_5_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_5
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_5_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_5_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_5_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_5_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_5_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_5
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_5_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_5_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_5_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_5_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_z(ccs_lp_piped_fp_mult_23_8_0_cmp_5_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_4_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_4_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_4_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_4_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_4_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_a;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_b;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_4_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_4_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_4_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_4_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_4_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_4_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_4_a_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_4_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_4_a_core
      = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_4_a_core[30:16]) , 16'b0000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_4_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_4_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_4_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_4_b_core
      = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_4_b_core[30:23]) , 23'b00000000000000000000000};
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_4 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_4_a),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_4_b),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_4_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_4_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_4_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_4_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_4_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_4_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_4_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_4_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_4
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_4_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_4_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_4_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_4_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_4_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_4
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_4_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_4_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_4_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_b_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_4_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_4_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_4_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_4_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_a(ccs_lp_piped_fp_mult_23_8_0_cmp_4_a),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_b(ccs_lp_piped_fp_mult_23_8_0_cmp_4_b),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_z(ccs_lp_piped_fp_mult_23_8_0_cmp_4_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_3
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_3 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_3_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_3_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_3_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_3_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_3_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_3_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_3_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_3_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_3_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_3_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_3_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_3_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_3_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_3_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_3_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_3_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_3 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_3_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_3_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_3_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_3_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_3_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_3_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_3_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_3_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_3_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_3_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_3_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_3
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_3_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_3_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_3_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_3_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_3_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_3_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_3_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_3
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_3_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_3_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_3_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_3_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_3_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_z(ccs_lp_piped_fp_mult_23_8_0_cmp_3_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_2_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_2_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_2_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_a;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_b;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_2_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_2_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_2_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_2_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_2_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_2_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_2_a_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_2_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_2_a_core
      = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_2_a_core[30:16]) , 16'b0000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_2_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_2_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_2_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_2_b_core
      = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_2_b_core[30:23]) , 23'b00000000000000000000000};
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_2 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_2_a),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_2_b),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_2_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_2_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_2_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_2_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_2_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_2_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_2_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_2_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_2
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_2_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_2_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_2_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_2
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_2_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_2_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_2_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_b_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_2_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_2_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_a(ccs_lp_piped_fp_mult_23_8_0_cmp_2_a),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_b(ccs_lp_piped_fp_mult_23_8_0_cmp_2_b),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_z(ccs_lp_piped_fp_mult_23_8_0_cmp_2_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_1_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_1_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_1_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_1_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_1_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_1_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_1_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_1_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_1 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_1_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_1_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_1_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_1_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_1_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_1_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_1_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_1_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_1_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_1_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_1
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_1_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_1_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_1
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_z(ccs_lp_piped_fp_mult_23_8_0_cmp_1_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_oswt_unreg, ccs_lp_piped_fp_mult_23_8_0_cmp_bawt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_a_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_b_core, ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_a;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_b;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_a_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_a_core
      = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_a_core[30:16]) , 16'b0000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_b_core
      = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_b_core[30:23]) , 23'b00000000000000000000000};
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_a),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_b),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp
      bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_b_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_a(ccs_lp_piped_fp_mult_23_8_0_cmp_a),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_b(ccs_lp_piped_fp_mult_23_8_0_cmp_b),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_z(ccs_lp_piped_fp_mult_23_8_0_cmp_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_11
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_11 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_11_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_11_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_11_a_core, ccs_lp_piped_fp_add_23_8_0_cmp_11_b_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_11_z_mxwt, ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_11_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_11_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_11_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_11_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_11_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_11_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_11_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_11_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_11_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_11_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_11_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_11_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_11_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_11_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_11_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp_11 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_11_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_11_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_11_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_11_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_11_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_11_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_11_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_11_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_11_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_11_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_11_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_11
      bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_11_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_11_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_11_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_11_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_11_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_11_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_11_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_11
      bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_11_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_11_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_11_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_11_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_11_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_11_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_z(ccs_lp_piped_fp_add_23_8_0_cmp_11_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_10
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_10 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_10_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_10_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_10_a_core, ccs_lp_piped_fp_add_23_8_0_cmp_10_b_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_10_z_mxwt, ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_10_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_10_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_10_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_10_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_10_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_10_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_10_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_10_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_10_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_10_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_10_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_10_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_10_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_10_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_10_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp_10 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_10_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_10_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_10_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_10_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_10_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_10_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_10_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_10_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_10_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_10_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_10_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_10
      bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_10_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_10_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_10_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_10_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_10_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_10_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_10_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_10
      bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_10_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_10_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_10_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_10_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_10_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_10_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_z(ccs_lp_piped_fp_add_23_8_0_cmp_10_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_9
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_9 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_9_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_9_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_9_a_core, ccs_lp_piped_fp_add_23_8_0_cmp_9_b_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_9_z_mxwt, ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_9_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_9_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_9_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_9_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_9_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_9_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_9_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_9_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_9_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_9_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_9_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_9_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_9_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_9_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_9_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp_9 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_9_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_9_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_9_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_9_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_9_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_9_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_9_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_9_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_9_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_9_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_9_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_9
      bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_9_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_9_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_9_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_9_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_9_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_9_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_9_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_9
      bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_9_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_9_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_9_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_9_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_9_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_9_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_z(ccs_lp_piped_fp_add_23_8_0_cmp_9_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_8
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_8 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_8_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_8_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_8_a_core, ccs_lp_piped_fp_add_23_8_0_cmp_8_b_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_8_z_mxwt, ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_8_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_8_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_8_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_8_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_8_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_8_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_8_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_8_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_8_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_8_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_8_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_8_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_8_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_8_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_8_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp_8 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_8_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_8_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_8_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_8_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_8_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_8_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_8_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_8_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_8_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_8_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_8_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_8
      bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_8_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_8_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_8_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_8_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_8_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_8_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_8_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_8
      bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_8_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_8_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_8_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_8_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_8_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_8_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_z(ccs_lp_piped_fp_add_23_8_0_cmp_8_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_7
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_7 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_7_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_7_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_7_a_core, ccs_lp_piped_fp_add_23_8_0_cmp_7_b_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_7_z_mxwt, ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_7_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_7_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_7_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_7_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_7_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_7_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_7_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_7_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_7_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_7_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_7_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_7_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_7_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_7_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_7_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp_7 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_7_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_7_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_7_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_7_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_7_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_7_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_7_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_7_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_7_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_7_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_7_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_7
      bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_7_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_7_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_7_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_7_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_7_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_7_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_7_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_7
      bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_7_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_7_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_7_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_7_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_7_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_7_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_z(ccs_lp_piped_fp_add_23_8_0_cmp_7_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_6
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_6 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_6_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_6_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_6_a_core, ccs_lp_piped_fp_add_23_8_0_cmp_6_b_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_6_z_mxwt, ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_6_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_6_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_6_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_6_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_6_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_6_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_6_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_6_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_6_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_6_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_6_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_6_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_6_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_6_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_6_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp_6 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_6_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_6_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_6_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_6_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_6_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_6_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_6_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_6_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_6_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_6_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_6_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_6
      bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_6_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_6_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_6_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_6_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_6_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_6_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_6_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_6
      bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_6_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_6_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_6_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_6_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_6_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_6_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_z(ccs_lp_piped_fp_add_23_8_0_cmp_6_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_5
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_5 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_5_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_5_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_5_a_core, ccs_lp_piped_fp_add_23_8_0_cmp_5_b_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_5_z_mxwt, ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_5_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_5_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_5_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_5_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_5_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_5_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_5_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_5_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_5_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_5_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_5_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_5_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_5_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_5_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_5_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp_5 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_5_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_5_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_5_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_5_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_5_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_5_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_5_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_5_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_5_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_5_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_5_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_5
      bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_5_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_5_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_5_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_5_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_5_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_5_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_5_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_5
      bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_5_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_5_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_5_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_5_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_5_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_5_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_z(ccs_lp_piped_fp_add_23_8_0_cmp_5_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_4
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_4 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_4_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_4_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_4_a_core, ccs_lp_piped_fp_add_23_8_0_cmp_4_b_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_4_z_mxwt, ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_4_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_4_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_4_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_4_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_4_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_4_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_4_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_4_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_4_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_4_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_4_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_4_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_4_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_4_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_4_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp_4 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_4_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_4_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_4_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_4_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_4_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_4_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_4_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_4_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_4_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_4_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_4_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_4
      bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_4_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_4_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_4_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_4_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_4_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_4_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_4_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_4
      bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_4_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_4_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_4_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_4_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_4_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_4_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_z(ccs_lp_piped_fp_add_23_8_0_cmp_4_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_3
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_3 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_3_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_3_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_3_a_core, ccs_lp_piped_fp_add_23_8_0_cmp_3_b_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_3_z_mxwt, ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_3_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_3_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_3_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_3_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_3_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_3_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_3_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_3_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_3_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_3_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_3_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_3_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_3_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_3_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_3_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp_3 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_3_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_3_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_3_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_3_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_3_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_3_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_3_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_3_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_3_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_3_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_3_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_3
      bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_3_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_3_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_3_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_3_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_3_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_3_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_3_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_3
      bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_3_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_3_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_3_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_3_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_3_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_3_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_z(ccs_lp_piped_fp_add_23_8_0_cmp_3_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_2
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_2 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_2_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_2_a_core, ccs_lp_piped_fp_add_23_8_0_cmp_2_b_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt, ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_2_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_2_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_2_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_2_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_2_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_2_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp_2 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_2_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_2_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_2_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_2_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_2_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_2_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_2_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_2_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_2_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_2_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_2
      bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_2_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_2_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_2_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_2
      bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_2_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_z(ccs_lp_piped_fp_add_23_8_0_cmp_2_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_1
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_1 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_1_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_1_a_core, ccs_lp_piped_fp_add_23_8_0_cmp_1_b_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt, ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_1_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_1_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_1_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_1_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_1_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_1_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp_1 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_1_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_1_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_1_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_1_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_1_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_1_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_1_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_1_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_1_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_1_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_1
      bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_1_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_1_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_1
      bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_z(ccs_lp_piped_fp_add_23_8_0_cmp_1_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp
// ------------------------------------------------------------------


module bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_oswt_unreg, ccs_lp_piped_fp_add_23_8_0_cmp_bawt,
      ccs_lp_piped_fp_add_23_8_0_cmp_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_a_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_b_core, ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_pipe_census)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl
      bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_iswt1_pff)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp
      bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_z(ccs_lp_piped_fp_add_23_8_0_cmp_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_bbox_resp_stream_rsci
// ------------------------------------------------------------------


module bbox_core_bbox_resp_stream_rsci (
  clk, arst_n, bbox_resp_stream_rsc_dat, bbox_resp_stream_rsc_vld, bbox_resp_stream_rsc_rdy,
      core_wen, bbox_resp_stream_rsci_oswt_unreg, bbox_resp_stream_rsci_bawt, bbox_resp_stream_rsci_iswt0,
      bbox_resp_stream_rsci_wen_comp, bbox_resp_stream_rsci_idat
);
  input clk;
  input arst_n;
  output [204:0] bbox_resp_stream_rsc_dat;
  output bbox_resp_stream_rsc_vld;
  input bbox_resp_stream_rsc_rdy;
  input core_wen;
  input bbox_resp_stream_rsci_oswt_unreg;
  output bbox_resp_stream_rsci_bawt;
  input bbox_resp_stream_rsci_iswt0;
  output bbox_resp_stream_rsci_wen_comp;
  input [204:0] bbox_resp_stream_rsci_idat;


  // Interconnect Declarations
  wire bbox_resp_stream_rsci_biwt;
  wire bbox_resp_stream_rsci_bdwt;
  wire bbox_resp_stream_rsci_bcwt;
  wire bbox_resp_stream_rsci_irdy;
  wire bbox_resp_stream_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd28),
  .width(32'sd205)) bbox_resp_stream_rsci (
      .irdy(bbox_resp_stream_rsci_irdy),
      .ivld(bbox_resp_stream_rsci_ivld_core_sct),
      .idat(bbox_resp_stream_rsci_idat),
      .rdy(bbox_resp_stream_rsc_rdy),
      .vld(bbox_resp_stream_rsc_vld),
      .dat(bbox_resp_stream_rsc_dat)
    );
  bbox_core_bbox_resp_stream_rsci_bbox_resp_stream_wait_ctrl bbox_core_bbox_resp_stream_rsci_bbox_resp_stream_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .bbox_resp_stream_rsci_oswt_unreg(bbox_resp_stream_rsci_oswt_unreg),
      .bbox_resp_stream_rsci_iswt0(bbox_resp_stream_rsci_iswt0),
      .bbox_resp_stream_rsci_biwt(bbox_resp_stream_rsci_biwt),
      .bbox_resp_stream_rsci_bdwt(bbox_resp_stream_rsci_bdwt),
      .bbox_resp_stream_rsci_bcwt(bbox_resp_stream_rsci_bcwt),
      .bbox_resp_stream_rsci_irdy(bbox_resp_stream_rsci_irdy),
      .bbox_resp_stream_rsci_ivld_core_sct(bbox_resp_stream_rsci_ivld_core_sct)
    );
  bbox_core_bbox_resp_stream_rsci_bbox_resp_stream_wait_dp bbox_core_bbox_resp_stream_rsci_bbox_resp_stream_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .bbox_resp_stream_rsci_oswt_unreg(bbox_resp_stream_rsci_oswt_unreg),
      .bbox_resp_stream_rsci_bawt(bbox_resp_stream_rsci_bawt),
      .bbox_resp_stream_rsci_wen_comp(bbox_resp_stream_rsci_wen_comp),
      .bbox_resp_stream_rsci_biwt(bbox_resp_stream_rsci_biwt),
      .bbox_resp_stream_rsci_bdwt(bbox_resp_stream_rsci_bdwt),
      .bbox_resp_stream_rsci_bcwt(bbox_resp_stream_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core_bbox_req_stream_rsci
// ------------------------------------------------------------------


module bbox_core_bbox_req_stream_rsci (
  clk, arst_n, bbox_req_stream_rsc_dat, bbox_req_stream_rsc_vld, bbox_req_stream_rsc_rdy,
      core_wen, bbox_req_stream_rsci_oswt_unreg, bbox_req_stream_rsci_bawt, bbox_req_stream_rsci_iswt0,
      bbox_req_stream_rsci_wen_comp, bbox_req_stream_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [385:0] bbox_req_stream_rsc_dat;
  input bbox_req_stream_rsc_vld;
  output bbox_req_stream_rsc_rdy;
  input core_wen;
  input bbox_req_stream_rsci_oswt_unreg;
  output bbox_req_stream_rsci_bawt;
  input bbox_req_stream_rsci_iswt0;
  output bbox_req_stream_rsci_wen_comp;
  output [385:0] bbox_req_stream_rsci_idat_mxwt;


  // Interconnect Declarations
  wire bbox_req_stream_rsci_biwt;
  wire bbox_req_stream_rsci_bdwt;
  wire bbox_req_stream_rsci_bcwt;
  wire bbox_req_stream_rsci_irdy_core_sct;
  wire bbox_req_stream_rsci_ivld;
  wire [385:0] bbox_req_stream_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd27),
  .width(32'sd386)) bbox_req_stream_rsci (
      .rdy(bbox_req_stream_rsc_rdy),
      .vld(bbox_req_stream_rsc_vld),
      .dat(bbox_req_stream_rsc_dat),
      .irdy(bbox_req_stream_rsci_irdy_core_sct),
      .ivld(bbox_req_stream_rsci_ivld),
      .idat(bbox_req_stream_rsci_idat)
    );
  bbox_core_bbox_req_stream_rsci_bbox_req_stream_wait_ctrl bbox_core_bbox_req_stream_rsci_bbox_req_stream_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .bbox_req_stream_rsci_oswt_unreg(bbox_req_stream_rsci_oswt_unreg),
      .bbox_req_stream_rsci_iswt0(bbox_req_stream_rsci_iswt0),
      .bbox_req_stream_rsci_biwt(bbox_req_stream_rsci_biwt),
      .bbox_req_stream_rsci_bdwt(bbox_req_stream_rsci_bdwt),
      .bbox_req_stream_rsci_bcwt(bbox_req_stream_rsci_bcwt),
      .bbox_req_stream_rsci_irdy_core_sct(bbox_req_stream_rsci_irdy_core_sct),
      .bbox_req_stream_rsci_ivld(bbox_req_stream_rsci_ivld)
    );
  bbox_core_bbox_req_stream_rsci_bbox_req_stream_wait_dp bbox_core_bbox_req_stream_rsci_bbox_req_stream_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .bbox_req_stream_rsci_oswt_unreg(bbox_req_stream_rsci_oswt_unreg),
      .bbox_req_stream_rsci_bawt(bbox_req_stream_rsci_bawt),
      .bbox_req_stream_rsci_wen_comp(bbox_req_stream_rsci_wen_comp),
      .bbox_req_stream_rsci_idat_mxwt(bbox_req_stream_rsci_idat_mxwt),
      .bbox_req_stream_rsci_biwt(bbox_req_stream_rsci_biwt),
      .bbox_req_stream_rsci_bdwt(bbox_req_stream_rsci_bdwt),
      .bbox_req_stream_rsci_bcwt(bbox_req_stream_rsci_bcwt),
      .bbox_req_stream_rsci_idat(bbox_req_stream_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_28
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_28 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_28_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_28_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_28_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_28_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_28_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_28_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_28_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_28_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_28_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_28_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_28_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_28_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_28_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_28_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_28_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_28_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_28_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_28_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_28_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_28_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_28_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_28_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_28_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_28_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_28 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_28_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_28_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_28_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_28_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_28_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_28_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_28_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_28_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_28_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_28_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_28_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_28
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_28_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_28_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_28_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_28_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_28_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_28_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_28_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_28_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_28_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_28_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_28_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_28_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_28_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_28_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_28_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_28
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_28_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_28_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_28_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_28_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_28_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_28_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_28_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_28_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_28_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_28_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_28_z(ccs_lp_piped_fp_mult_23_8_0_cmp_28_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_27
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_27 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_27_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_27_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_27_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_27_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_27_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_27_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_27_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_27_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_27_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_27_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_27_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_27_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_27_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_27_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_27_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_27_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_27_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_27_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_27_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_27_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_27_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_27_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_27_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_27_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_27 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_27_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_27_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_27_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_27_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_27_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_27_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_27_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_27_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_27_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_27_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_27_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_27
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_27_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_27_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_27_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_27_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_27_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_27_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_27_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_27_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_27_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_27_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_27_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_27_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_27_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_27_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_27_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_27
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_27_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_27_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_27_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_27_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_27_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_27_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_27_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_27_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_27_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_27_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_27_z(ccs_lp_piped_fp_mult_23_8_0_cmp_27_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_26
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_26 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_26_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_26_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_26_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_26_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_26_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_26_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_26_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_26_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_26_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_26_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_26_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_26_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_26_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_26_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_26_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_26_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_26_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_26_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_26_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_26_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_26_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_26_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_26_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_26_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_26 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_26_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_26_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_26_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_26_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_26_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_26_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_26_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_26_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_26_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_26_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_26_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_26
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_26_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_26_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_26_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_26_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_26_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_26_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_26_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_26_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_26_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_26_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_26_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_26_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_26_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_26_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_26_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_26
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_26_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_26_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_26_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_26_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_26_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_26_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_26_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_26_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_26_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_26_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_26_z(ccs_lp_piped_fp_mult_23_8_0_cmp_26_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_25
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_25 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_25_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_25_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_25_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_25_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_25_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_25_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_25_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_25_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_25_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_25_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_25_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_25_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_25_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_25_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_25_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_25_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_25_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_25_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_25_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_25_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_25_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_25_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_25_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_25_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_25 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_25_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_25_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_25_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_25_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_25_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_25_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_25_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_25_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_25_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_25_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_25_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_25
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_25_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_25_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_25_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_25_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_25_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_25_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_25_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_25_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_25_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_25_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_25_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_25_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_25_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_25_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_25_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_25
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_25_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_25_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_25_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_25_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_25_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_25_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_25_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_25_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_25_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_25_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_25_z(ccs_lp_piped_fp_mult_23_8_0_cmp_25_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_24
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_24 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_24_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_24_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_24_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_24_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_24_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_24_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_24_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_24_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_24_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_24_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_24_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_24_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_24_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_24_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_24_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_24_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_24_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_24_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_24_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_24_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_24_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_24_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_24_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_24_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_24 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_24_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_24_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_24_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_24_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_24_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_24_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_24_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_24_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_24_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_24_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_24_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_24
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_24_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_24_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_24_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_24_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_24_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_24_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_24_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_24_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_24_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_24_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_24_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_24_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_24_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_24_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_24_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_24
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_24_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_24_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_24_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_24_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_24_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_24_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_24_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_24_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_24_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_24_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_24_z(ccs_lp_piped_fp_mult_23_8_0_cmp_24_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_23
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_23 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_23_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_23_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_23_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_23_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_23_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_23_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_23_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_23_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_23_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_23_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_23_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_23_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_23_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_23_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_23 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_23_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_23_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_23_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_23_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_23_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_23_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_23_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_23_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_23_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_23_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_23_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_23
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_23_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_23_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_23_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_23_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_23_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_23_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_23
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_23_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_23_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_23_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_23_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_23_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_z(ccs_lp_piped_fp_mult_23_8_0_cmp_23_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_22_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_22_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_22_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_22_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_22_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_22_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_22_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_22_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_22_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_22_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_22_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_22 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_22_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_22_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_22_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_22_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_22_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_22_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_22_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_22_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_22_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_22_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_22
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_22_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_22_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_22_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_22_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_22_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_22
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_22_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_22_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_22_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_22_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_z(ccs_lp_piped_fp_mult_23_8_0_cmp_22_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_21
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_21 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_21_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_21_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_21_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_21_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_21_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_21_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_21_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_21_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_21_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_21_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_21_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_21_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_21_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_21_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_21_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_21_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_21 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_21_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_21_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_21_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_21_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_21_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_21_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_21_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_21_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_21_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_21_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_21_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_21
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_21_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_21_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_21_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_21_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_21_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_21_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_21_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_21
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_21_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_21_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_21_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_21_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_21_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_z(ccs_lp_piped_fp_mult_23_8_0_cmp_21_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_20_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_20_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_20_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_20_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_20_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_20_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_20_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_20_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_20_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_20_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_20_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_20 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_20_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_20_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_20_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_20_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_20_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_20_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_20_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_20_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_20_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_20_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_20
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_20_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_20_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_20_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_20_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_20_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_20
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_20_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_20_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_20_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_20_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_z(ccs_lp_piped_fp_mult_23_8_0_cmp_20_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_19
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_19 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_19_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_19_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_19_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_19_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_19_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_19_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_19_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_19_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_19_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_19_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_19_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_19_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_19_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_19_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_19_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_19_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_19 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_19_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_19_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_19_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_19_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_19_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_19_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_19_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_19_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_19_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_19_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_19_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_19
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_19_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_19_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_19_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_19_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_19_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_19_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_19_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_19
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_19_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_19_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_19_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_19_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_19_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_z(ccs_lp_piped_fp_mult_23_8_0_cmp_19_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_18_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_18_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_18_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_18_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_18_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_18_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_18_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_18_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_18_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_18_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_18_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_18 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_18_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_18_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_18_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_18_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_18_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_18_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_18_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_18_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_18_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_18_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_18
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_18_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_18_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_18_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_18_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_18_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_18
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_18_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_18_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_18_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_18_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_z(ccs_lp_piped_fp_mult_23_8_0_cmp_18_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_17
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_17 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_17_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_17_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_17_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_17_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_17_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_17_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_17_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_17_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_17_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_17_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_17_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_17_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_17_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_17_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_17_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_17_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_17 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_17_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_17_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_17_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_17_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_17_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_17_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_17_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_17_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_17_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_17_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_17_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_17
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_17_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_17_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_17_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_17_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_17_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_17_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_17_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_17
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_17_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_17_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_17_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_17_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_17_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_z(ccs_lp_piped_fp_mult_23_8_0_cmp_17_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_16_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_16_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_16_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_16_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_16_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_16_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_16_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_16_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_16_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_16_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_16_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_16 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_16_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_16_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_16_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_16_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_16_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_16_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_16_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_16_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_16_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_16_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_16
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_16_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_16_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_16_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_16_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_16_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_16
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_16_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_16_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_16_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_16_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_z(ccs_lp_piped_fp_mult_23_8_0_cmp_16_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_15
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_15 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_15_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_15_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_15_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_15_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_15_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_15_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_15_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_15_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_15_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_15_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_15_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_15_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_15_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_15_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_15_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_15_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_15 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_15_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_15_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_15_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_15_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_15_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_15_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_15_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_15_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_15_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_15_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_15_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_15
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_15_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_15_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_15_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_15_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_15_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_15_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_15_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_15
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_15_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_15_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_15_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_15_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_15_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_z(ccs_lp_piped_fp_mult_23_8_0_cmp_15_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_14_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_14_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_14_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_14_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_14_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_14_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_14_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_14_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_14_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_14_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_14_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_14 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_14_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_14_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_14_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_14_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_14_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_14_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_14_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_14_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_14_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_14_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_14
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_14_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_14_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_14_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_14_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_14_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_14
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_14_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_14_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_14_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_14_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_z(ccs_lp_piped_fp_mult_23_8_0_cmp_14_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_13
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_13 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_13_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_13_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_13_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_13_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_13_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_13_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_13_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_13_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_13_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_13_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_13_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_13_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_13_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_13_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_13_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_13_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_13 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_13_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_13_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_13_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_13_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_13_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_13_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_13_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_13_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_13_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_13_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_13_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_13
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_13_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_13_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_13_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_13_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_13_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_13_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_13_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_13
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_13_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_13_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_13_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_13_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_13_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_z(ccs_lp_piped_fp_mult_23_8_0_cmp_13_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_12_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_12_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_12_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_12_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_12_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_12_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_12_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_12_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_12_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_12_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_12_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_12 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_12_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_12_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_12_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_12_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_12_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_12_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_12_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_12_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_12_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_12_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_12
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_12_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_12_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_12_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_12_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_12_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_12
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_12_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_12_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_12_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_12_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_z(ccs_lp_piped_fp_mult_23_8_0_cmp_12_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_11
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_11 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_11_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_11_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_11_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_11_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_11_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_11_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_11_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_11_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_11_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_11_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_11_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_11_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_11_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_11_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_11_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_11_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_11 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_11_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_11_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_11_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_11_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_11_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_11_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_11_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_11_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_11_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_11_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_11_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_11
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_11_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_11_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_11_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_11_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_11_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_11_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_11_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_11
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_11_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_11_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_11_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_11_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_11_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_z(ccs_lp_piped_fp_mult_23_8_0_cmp_11_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_10_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_10_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_10_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_10_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_10_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_10_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_10_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_10_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_10_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_10_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_10_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_10 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_10_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_10_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_10_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_10_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_10_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_10_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_10_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_10_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_10_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_10_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_10
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_10_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_10_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_10_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_10_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_10_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_10
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_10_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_10_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_10_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_10_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_z(ccs_lp_piped_fp_mult_23_8_0_cmp_10_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_9
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_9 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_9_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_9_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_9_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_9_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_9_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_9_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_9_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_9_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_9_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_9_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_9_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_9_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_9_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_9_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_9_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_9_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_9 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_9_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_9_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_9_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_9_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_9_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_9_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_9_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_9_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_9_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_9_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_9_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_9
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_9_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_9_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_9_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_9_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_9_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_9_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_9_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_9
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_9_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_9_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_9_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_9_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_9_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_z(ccs_lp_piped_fp_mult_23_8_0_cmp_9_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_8_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_8_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_8_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_8_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_8_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_8_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_8_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_8_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_8_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_8_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_8_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_8 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_8_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_8_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_8_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_8_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_8_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_8_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_8_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_8_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_8_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_8_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_8
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_8_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_8_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_8_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_8_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_8_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_8
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_8_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_8_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_8_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_8_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_z(ccs_lp_piped_fp_mult_23_8_0_cmp_8_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_7
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_7 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_7_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_7_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_7_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_7_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_7_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_7_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_7_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_7_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_7_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_7_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_7_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_7_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_7_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_7_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_7_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_7_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_7 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_7_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_7_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_7_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_7_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_7_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_7_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_7_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_7_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_7_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_7_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_7_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_7
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_7_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_7_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_7_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_7_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_7_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_7_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_7_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_7
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_7_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_7_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_7_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_7_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_7_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_z(ccs_lp_piped_fp_mult_23_8_0_cmp_7_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_6_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_6_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_6_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_6_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_6_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_6_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_6_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_6_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_6_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_6_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_6_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_6 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_6_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_6_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_6_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_6_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_6_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_6_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_6_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_6_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_6_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_6_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_6
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_6_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_6_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_6_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_6_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_6_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_6
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_6_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_6_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_6_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_6_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_z(ccs_lp_piped_fp_mult_23_8_0_cmp_6_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_5_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_5_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_5_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_5_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_5_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_5_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_5_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_5_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_5_a;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_5_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_5_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_5_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_5_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_5_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_5_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_5_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_5_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_5_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_5_a_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_5_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_5_a_core
      = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_5_a_core[30:0])};
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_5 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_5_a),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_5_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_5_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_5_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_5_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_5_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_5_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_5_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_5_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_5_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_5
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_5_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_5_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_5_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_5_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_5_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_5
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_5_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_5_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_a_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_5_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_5_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_5_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_5_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_a(ccs_lp_piped_fp_mult_23_8_0_cmp_5_a),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_z(ccs_lp_piped_fp_mult_23_8_0_cmp_5_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_4_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_4_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_4_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_4_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_4_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_a;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_4_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_4_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_4_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_4_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_4_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_4_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_4_a_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_4_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_4_a_core
      = {1'b0 , (ccs_lp_piped_fp_mult_23_8_0_cmp_4_a_core[30:0])};
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_4 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_4_a),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_4_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_4_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_4_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_4_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_4_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_4_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_4_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_4_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_4_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_4
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_4_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_4_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_4_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_4_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_4_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_4
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_4_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_a_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_4_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_4_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_4_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_4_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_a(ccs_lp_piped_fp_mult_23_8_0_cmp_4_a),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_z(ccs_lp_piped_fp_mult_23_8_0_cmp_4_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_3
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_3 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_3_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_3_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_3_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_3_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_3_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_3_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_3_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_3_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_3_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_3_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_3_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_3_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_3_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_3_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_3_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_3_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_3 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_3_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_3_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_3_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_3_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_3_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_3_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_3_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_3_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_3_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_3_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_3_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_3
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_3_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_3_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_3_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_3_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_3_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_3_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_3_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_3
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_3_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_3_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_3_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_3_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_3_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_z(ccs_lp_piped_fp_mult_23_8_0_cmp_3_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_2_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_2_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_2_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_2_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_2_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_2_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_2_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_2_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_2 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_2_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_2_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_2_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_2_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_2_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_2_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_2_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_2_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_2_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_2_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_2
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_2_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_2_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_2_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_2
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_2_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_2_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_2_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_z(ccs_lp_piped_fp_mult_23_8_0_cmp_2_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_1_oswt_unreg,
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt, ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1,
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_a_core, ccs_lp_piped_fp_mult_23_8_0_cmp_1_b_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt, ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_1_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_1_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_1_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_1_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_1_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_1_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp_1 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_1_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_1_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_1_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_1_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_1_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_1_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_1_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_1_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_1_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_1_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_1
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_1_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_1_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_1
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_1_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_1_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_z(ccs_lp_piped_fp_mult_23_8_0_cmp_1_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_mult_23_8_0_cmp_oswt_unreg, ccs_lp_piped_fp_mult_23_8_0_cmp_bawt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1, ccs_lp_piped_fp_mult_23_8_0_cmp_a_core,
      ccs_lp_piped_fp_mult_23_8_0_cmp_b_core, ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt,
      ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_oswt_unreg;
  output ccs_lp_piped_fp_mult_23_8_0_cmp_bawt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_a_core;
  input [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_b_core;
  output [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt;
  input ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_biwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_z;
  wire [7:0] ccs_lp_piped_fp_mult_23_8_0_cmp_status;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_launch_core_sct;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_pipe_full;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_pipe_ovf;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_arrive;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_push_out_n;
  wire [1:0] ccs_lp_piped_fp_mult_23_8_0_cmp_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_mult_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_mult_23_8_0_cmp (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_mult_23_8_0_cmp_a_core),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_mult_23_8_0_cmp_z),
      .status(ccs_lp_piped_fp_mult_23_8_0_cmp_status),
      .launch(ccs_lp_piped_fp_mult_23_8_0_cmp_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_mult_23_8_0_cmp_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_mult_23_8_0_cmp_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_mult_23_8_0_cmp_arrive),
      .push_out_n(ccs_lp_piped_fp_mult_23_8_0_cmp_push_out_n),
      .pipe_census(ccs_lp_piped_fp_mult_23_8_0_cmp_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_oswt_unreg(ccs_lp_piped_fp_mult_23_8_0_cmp_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_launch_core_sct(ccs_lp_piped_fp_mult_23_8_0_cmp_launch_core_sct),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1_pff(ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp
      ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_ccs_dw_lp_piped_fp_mult_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_biwt(ccs_lp_piped_fp_mult_23_8_0_cmp_biwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt(ccs_lp_piped_fp_mult_23_8_0_cmp_bdwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_z(ccs_lp_piped_fp_mult_23_8_0_cmp_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_17
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_17 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_17_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_17_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_17_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_17_a_core, ccs_lp_piped_fp_add_23_8_0_cmp_17_b_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_17_z_mxwt, ccs_lp_piped_fp_add_23_8_0_cmp_17_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_17_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_17_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_17_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_17_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_17_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_17_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_17_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_17_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_17_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_17_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_17_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_17_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_17_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_17_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_17_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_17_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_17_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp_17 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_17_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_17_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_17_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_17_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_17_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_17_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_17_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_17_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_17_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_17_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_17_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_17
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_17_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_17_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_17_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_17_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_17_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_17_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_17_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_17_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_17_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_17_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_17_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_17_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_17_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_17_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_17_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_17
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_17_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_17_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_17_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_17_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_17_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_17_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_17_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_17_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_17_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_17_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_17_z(ccs_lp_piped_fp_add_23_8_0_cmp_17_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_16
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_16 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_16_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_16_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_16_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_16_a_core, ccs_lp_piped_fp_add_23_8_0_cmp_16_b_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_16_z_mxwt, ccs_lp_piped_fp_add_23_8_0_cmp_16_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_16_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_16_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_16_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_16_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_16_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_16_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_16_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_16_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_16_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_16_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_16_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_16_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_16_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_16_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_16_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_16_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_16_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp_16 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_16_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_16_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_16_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_16_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_16_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_16_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_16_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_16_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_16_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_16_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_16_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_16
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_16_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_16_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_16_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_16_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_16_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_16_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_16_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_16_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_16_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_16_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_16_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_16_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_16_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_16_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_16_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_16
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_16_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_16_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_16_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_16_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_16_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_16_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_16_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_16_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_16_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_16_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_16_z(ccs_lp_piped_fp_add_23_8_0_cmp_16_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_15
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_15 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_15_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_15_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_15_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_15_a_core, ccs_lp_piped_fp_add_23_8_0_cmp_15_b_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_15_z_mxwt, ccs_lp_piped_fp_add_23_8_0_cmp_15_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_15_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_15_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_15_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_15_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_15_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_15_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_15_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_15_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_15_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_15_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_15_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_15_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_15_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_15_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_15_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_15_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_15_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp_15 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_15_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_15_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_15_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_15_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_15_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_15_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_15_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_15_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_15_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_15_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_15_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_15
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_15_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_15_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_15_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_15_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_15_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_15_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_15_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_15_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_15_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_15_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_15_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_15_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_15_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_15_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_15_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_15
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_15_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_15_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_15_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_15_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_15_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_15_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_15_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_15_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_15_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_15_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_15_z(ccs_lp_piped_fp_add_23_8_0_cmp_15_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_14
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_14 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_14_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_14_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_14_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_14_a_core, ccs_lp_piped_fp_add_23_8_0_cmp_14_b_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_14_z_mxwt, ccs_lp_piped_fp_add_23_8_0_cmp_14_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_14_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_14_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_14_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_14_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_14_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_14_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_14_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_14_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_14_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_14_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_14_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_14_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_14_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_14_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_14_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_14_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_14_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp_14 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_14_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_14_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_14_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_14_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_14_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_14_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_14_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_14_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_14_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_14_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_14_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_14
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_14_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_14_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_14_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_14_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_14_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_14_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_14_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_14_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_14_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_14_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_14_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_14_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_14_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_14_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_14_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_14
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_14_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_14_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_14_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_14_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_14_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_14_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_14_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_14_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_14_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_14_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_14_z(ccs_lp_piped_fp_add_23_8_0_cmp_14_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_13
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_13 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_13_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_13_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_13_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_13_a_core, ccs_lp_piped_fp_add_23_8_0_cmp_13_b_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_13_z_mxwt, ccs_lp_piped_fp_add_23_8_0_cmp_13_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_13_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_13_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_13_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_13_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_13_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_13_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_13_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_13_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_13_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_13_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_13_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_13_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_13_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_13_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_13_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_13_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_13_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp_13 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_13_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_13_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_13_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_13_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_13_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_13_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_13_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_13_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_13_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_13_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_13_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_13
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_13_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_13_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_13_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_13_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_13_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_13_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_13_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_13_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_13_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_13_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_13_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_13_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_13_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_13_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_13_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_13
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_13_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_13_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_13_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_13_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_13_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_13_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_13_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_13_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_13_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_13_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_13_z(ccs_lp_piped_fp_add_23_8_0_cmp_13_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_12
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_12 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_12_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_12_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_12_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_12_a_core, ccs_lp_piped_fp_add_23_8_0_cmp_12_b_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_12_z_mxwt, ccs_lp_piped_fp_add_23_8_0_cmp_12_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_12_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_12_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_12_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_12_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_12_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_12_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_12_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_12_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_12_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_12_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_12_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_12_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_12_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_12_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_12_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_12_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_12_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp_12 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_12_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_12_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_12_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_12_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_12_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_12_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_12_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_12_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_12_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_12_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_12_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_12
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_12_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_12_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_12_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_12_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_12_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_12_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_12_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_12_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_12_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_12_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_12_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_12_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_12_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_12_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_12_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_12
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_12_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_12_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_12_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_12_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_12_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_12_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_12_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_12_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_12_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_12_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_12_z(ccs_lp_piped_fp_add_23_8_0_cmp_12_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_11
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_11 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_11_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_11_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_11_a_core, ccs_lp_piped_fp_add_23_8_0_cmp_11_b_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_11_z_mxwt, ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_11_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_11_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_11_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_11_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_11_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_11_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_11_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_11_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_11_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_11_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_11_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_11_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_11_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_11_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_11_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp_11 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_11_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_11_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_11_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_11_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_11_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_11_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_11_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_11_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_11_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_11_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_11_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_11
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_11_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_11_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_11_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_11_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_11_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_11_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_11_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_11
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_11_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_11_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_11_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_11_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_11_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_11_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_z(ccs_lp_piped_fp_add_23_8_0_cmp_11_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_10
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_10 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_10_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_10_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_10_a_core, ccs_lp_piped_fp_add_23_8_0_cmp_10_b_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_10_z_mxwt, ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_10_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_10_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_10_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_10_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_10_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_10_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_10_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_10_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_10_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_10_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_10_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_10_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_10_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_10_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_10_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp_10 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_10_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_10_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_10_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_10_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_10_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_10_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_10_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_10_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_10_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_10_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_10_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_10
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_10_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_10_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_10_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_10_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_10_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_10_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_10_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_10
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_10_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_10_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_10_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_10_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_10_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_10_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_z(ccs_lp_piped_fp_add_23_8_0_cmp_10_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_9
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_9 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_9_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_9_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_9_a_core, ccs_lp_piped_fp_add_23_8_0_cmp_9_b_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_9_z_mxwt, ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_9_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_9_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_9_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_9_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_9_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_9_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_9_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_9_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_9_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_9_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_9_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_9_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_9_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_9_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_9_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp_9 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_9_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_9_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_9_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_9_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_9_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_9_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_9_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_9_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_9_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_9_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_9_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_9
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_9_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_9_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_9_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_9_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_9_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_9_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_9_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_9
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_9_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_9_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_9_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_9_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_9_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_9_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_z(ccs_lp_piped_fp_add_23_8_0_cmp_9_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_8
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_8 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_8_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_8_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_8_a_core, ccs_lp_piped_fp_add_23_8_0_cmp_8_b_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_8_z_mxwt, ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_8_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_8_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_8_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_8_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_8_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_8_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_8_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_8_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_8_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_8_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_8_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_8_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_8_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_8_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_8_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp_8 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_8_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_8_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_8_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_8_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_8_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_8_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_8_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_8_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_8_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_8_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_8_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_8
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_8_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_8_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_8_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_8_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_8_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_8_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_8_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_8
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_8_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_8_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_8_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_8_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_8_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_8_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_z(ccs_lp_piped_fp_add_23_8_0_cmp_8_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_7
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_7 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_7_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_7_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_7_a_core, ccs_lp_piped_fp_add_23_8_0_cmp_7_b_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_7_z_mxwt, ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_7_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_7_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_7_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_7_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_7_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_7_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_7_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_7_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_7_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_7_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_7_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_7_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_7_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_7_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_7_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp_7 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_7_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_7_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_7_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_7_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_7_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_7_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_7_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_7_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_7_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_7_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_7_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_7
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_7_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_7_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_7_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_7_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_7_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_7_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_7_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_7
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_7_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_7_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_7_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_7_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_7_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_7_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_z(ccs_lp_piped_fp_add_23_8_0_cmp_7_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_6
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_6 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_6_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_6_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_6_a_core, ccs_lp_piped_fp_add_23_8_0_cmp_6_b_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_6_z_mxwt, ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_6_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_6_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_6_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_6_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_6_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_6_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_6_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_6_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_6_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_6_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_6_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_6_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_6_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_6_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_6_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp_6 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_6_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_6_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_6_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_6_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_6_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_6_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_6_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_6_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_6_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_6_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_6_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_6
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_6_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_6_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_6_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_6_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_6_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_6_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_6_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_6
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_6_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_6_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_6_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_6_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_6_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_6_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_z(ccs_lp_piped_fp_add_23_8_0_cmp_6_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_5
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_5 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_5_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_5_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_5_a_core, ccs_lp_piped_fp_add_23_8_0_cmp_5_b_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_5_z_mxwt, ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_5_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_5_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_5_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_5_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_5_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_5_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_5_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_5_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_5_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_5_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_5_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_5_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_5_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_5_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_5_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp_5 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_5_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_5_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_5_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_5_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_5_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_5_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_5_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_5_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_5_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_5_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_5_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_5
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_5_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_5_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_5_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_5_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_5_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_5_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_5_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_5
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_5_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_5_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_5_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_5_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_5_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_5_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_z(ccs_lp_piped_fp_add_23_8_0_cmp_5_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_4
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_4 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_4_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_4_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_4_a_core, ccs_lp_piped_fp_add_23_8_0_cmp_4_b_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_4_z_mxwt, ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_4_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_4_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_4_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_4_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_4_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_4_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_4_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_4_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_4_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_4_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_4_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_4_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_4_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_4_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_4_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp_4 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_4_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_4_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_4_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_4_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_4_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_4_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_4_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_4_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_4_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_4_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_4_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_4
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_4_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_4_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_4_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_4_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_4_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_4_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_4_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_4
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_4_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_4_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_4_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_4_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_4_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_4_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_z(ccs_lp_piped_fp_add_23_8_0_cmp_4_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_3
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_3 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_3_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_3_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_3_a_core, ccs_lp_piped_fp_add_23_8_0_cmp_3_b_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_3_z_mxwt, ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_3_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_3_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_3_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_3_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_3_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_3_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_3_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_3_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_3_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_3_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_3_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_3_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_3_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_3_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_3_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp_3 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_3_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_3_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_3_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_3_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_3_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_3_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_3_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_3_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_3_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_3_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_3_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_3
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_3_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_3_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_3_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_3_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_3_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_3_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_3_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_3
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_3_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_3_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_3_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_3_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_3_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_3_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_z(ccs_lp_piped_fp_add_23_8_0_cmp_3_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_2
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_2 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_2_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_2_a_core, ccs_lp_piped_fp_add_23_8_0_cmp_2_b_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt, ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_2_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_2_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_2_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_2_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_2_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_2_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp_2 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_2_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_2_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_2_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_2_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_2_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_2_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_2_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_2_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_2_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_2_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_2
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_2_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_2_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_2_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_2
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_2_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_2_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_2_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_z(ccs_lp_piped_fp_add_23_8_0_cmp_2_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_1
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_1 (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_1_oswt_unreg,
      ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt, ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1,
      ccs_lp_piped_fp_add_23_8_0_cmp_1_a_core, ccs_lp_piped_fp_add_23_8_0_cmp_1_b_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt, ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_1_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_1_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_1_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_1_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_1_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_1_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp_1 (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_1_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_1_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_1_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_1_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_1_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_1_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_1_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_1_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_1_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_1_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_1
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_1_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_1_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_1
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_1_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_1_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_z(ccs_lp_piped_fp_add_23_8_0_cmp_1_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_add_23_8_0_cmp
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_add_23_8_0_cmp (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_add_23_8_0_cmp_oswt_unreg, ccs_lp_piped_fp_add_23_8_0_cmp_bawt,
      ccs_lp_piped_fp_add_23_8_0_cmp_iswt1, ccs_lp_piped_fp_add_23_8_0_cmp_a_core,
      ccs_lp_piped_fp_add_23_8_0_cmp_b_core, ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_add_23_8_0_cmp_oswt_unreg;
  output ccs_lp_piped_fp_add_23_8_0_cmp_bawt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_iswt1;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_a_core;
  input [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_b_core;
  output [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt;
  input ccs_lp_piped_fp_add_23_8_0_cmp_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_add_23_8_0_cmp_biwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_bdwt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_z;
  wire [7:0] ccs_lp_piped_fp_add_23_8_0_cmp_status;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_launch_core_sct;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_pipe_full;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_pipe_ovf;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_arrive;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_push_out_n;
  wire [1:0] ccs_lp_piped_fp_add_23_8_0_cmp_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  ccs_dw_lp_piped_fp_add_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_add_23_8_0_cmp (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_a_core),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_b_core),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_add_23_8_0_cmp_z),
      .status(ccs_lp_piped_fp_add_23_8_0_cmp_status),
      .launch(ccs_lp_piped_fp_add_23_8_0_cmp_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_add_23_8_0_cmp_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_add_23_8_0_cmp_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_add_23_8_0_cmp_arrive),
      .push_out_n(ccs_lp_piped_fp_add_23_8_0_cmp_push_out_n),
      .pipe_census(ccs_lp_piped_fp_add_23_8_0_cmp_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_ctrl_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_oswt_unreg(ccs_lp_piped_fp_add_23_8_0_cmp_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_launch_core_sct(ccs_lp_piped_fp_add_23_8_0_cmp_launch_core_sct),
      .ccs_lp_piped_fp_add_23_8_0_cmp_iswt1_pff(ccs_lp_piped_fp_add_23_8_0_cmp_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp
      ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_ccs_dw_lp_piped_fp_add_23_8_0_1_2_0_0_1_0_0_0_4_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_add_23_8_0_cmp_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_biwt(ccs_lp_piped_fp_add_23_8_0_cmp_biwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_bdwt(ccs_lp_piped_fp_add_23_8_0_cmp_bdwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_z(ccs_lp_piped_fp_add_23_8_0_cmp_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ccs_lp_piped_fp_recip_23_8_0_cmp
// ------------------------------------------------------------------


module ist_core_ccs_lp_piped_fp_recip_23_8_0_cmp (
  clk, arst_n, core_wen, core_wten, ccs_lp_piped_fp_recip_23_8_0_cmp_oswt_unreg,
      ccs_lp_piped_fp_recip_23_8_0_cmp_bawt, ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1,
      ccs_lp_piped_fp_recip_23_8_0_cmp_a_core, ccs_lp_piped_fp_recip_23_8_0_cmp_z_mxwt,
      ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1_pff
);
  input clk;
  input arst_n;
  input core_wen;
  input core_wten;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_oswt_unreg;
  output ccs_lp_piped_fp_recip_23_8_0_cmp_bawt;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1;
  input [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_a_core;
  output [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_z_mxwt;
  input ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1_pff;


  // Interconnect Declarations
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_biwt;
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_bdwt;
  wire [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_a;
  wire [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_z;
  wire [7:0] ccs_lp_piped_fp_recip_23_8_0_cmp_status;
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_launch_core_sct;
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_pipe_full;
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_pipe_ovf;
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_arrive;
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_push_out_n;
  wire [1:0] ccs_lp_piped_fp_recip_23_8_0_cmp_pipe_census;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_recip_23_8_0_cmp_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_dp_inst_ccs_lp_piped_fp_recip_23_8_0_cmp_a_core;
  assign nl_ist_core_ccs_lp_piped_fp_recip_23_8_0_cmp_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_dp_inst_ccs_lp_piped_fp_recip_23_8_0_cmp_a_core
      = {1'b0 , (ccs_lp_piped_fp_recip_23_8_0_cmp_a_core[30:0])};
  ccs_dw_lp_piped_fp_recip_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0),
  .in_reg(32'sd1),
  .stages(32'sd2),
  .out_reg(32'sd0),
  .no_pm(32'sd0),
  .has_rst_a(32'sd1),
  .has_rst_s(32'sd0),
  .ph_arst(32'sd0),
  .ph_srst(32'sd0)) ccs_lp_piped_fp_recip_23_8_0_cmp (
      .clk(clk),
      .a_rst(arst_n),
      .s_rst(1'b1),
      .a(ccs_lp_piped_fp_recip_23_8_0_cmp_a),
      .rnd(3'b000),
      .z(ccs_lp_piped_fp_recip_23_8_0_cmp_z),
      .status(ccs_lp_piped_fp_recip_23_8_0_cmp_status),
      .launch(ccs_lp_piped_fp_recip_23_8_0_cmp_launch_core_sct),
      .pipe_full(ccs_lp_piped_fp_recip_23_8_0_cmp_pipe_full),
      .pipe_ovf(ccs_lp_piped_fp_recip_23_8_0_cmp_pipe_ovf),
      .accept_n(1'b0),
      .arrive(ccs_lp_piped_fp_recip_23_8_0_cmp_arrive),
      .push_out_n(ccs_lp_piped_fp_recip_23_8_0_cmp_push_out_n),
      .pipe_census(ccs_lp_piped_fp_recip_23_8_0_cmp_pipe_census)
    );
  ist_core_ccs_lp_piped_fp_recip_23_8_0_cmp_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_ctrl
      ist_core_ccs_lp_piped_fp_recip_23_8_0_cmp_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_ctrl_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_oswt_unreg(ccs_lp_piped_fp_recip_23_8_0_cmp_oswt_unreg),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1(ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_biwt(ccs_lp_piped_fp_recip_23_8_0_cmp_biwt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_bdwt(ccs_lp_piped_fp_recip_23_8_0_cmp_bdwt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_launch_core_sct(ccs_lp_piped_fp_recip_23_8_0_cmp_launch_core_sct),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1_pff(ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1_pff)
    );
  ist_core_ccs_lp_piped_fp_recip_23_8_0_cmp_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_dp
      ist_core_ccs_lp_piped_fp_recip_23_8_0_cmp_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_bawt(ccs_lp_piped_fp_recip_23_8_0_cmp_bawt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_a_core(nl_ist_core_ccs_lp_piped_fp_recip_23_8_0_cmp_ccs_dw_lp_piped_fp_recip_23_8_0_1_2_0_0_1_0_0_0_2_wait_dp_inst_ccs_lp_piped_fp_recip_23_8_0_cmp_a_core[31:0]),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_z_mxwt(ccs_lp_piped_fp_recip_23_8_0_cmp_z_mxwt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_biwt(ccs_lp_piped_fp_recip_23_8_0_cmp_biwt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_bdwt(ccs_lp_piped_fp_recip_23_8_0_cmp_bdwt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_a(ccs_lp_piped_fp_recip_23_8_0_cmp_a),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_z(ccs_lp_piped_fp_recip_23_8_0_cmp_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ist_resp_stream_rsci
// ------------------------------------------------------------------


module ist_core_ist_resp_stream_rsci (
  clk, arst_n, ist_resp_stream_rsc_dat, ist_resp_stream_rsc_vld, ist_resp_stream_rsc_rdy,
      core_wen, ist_resp_stream_rsci_oswt_unreg, ist_resp_stream_rsci_bawt, ist_resp_stream_rsci_iswt0,
      ist_resp_stream_rsci_wen_comp, ist_resp_stream_rsci_idat
);
  input clk;
  input arst_n;
  output [106:0] ist_resp_stream_rsc_dat;
  output ist_resp_stream_rsc_vld;
  input ist_resp_stream_rsc_rdy;
  input core_wen;
  input ist_resp_stream_rsci_oswt_unreg;
  output ist_resp_stream_rsci_bawt;
  input ist_resp_stream_rsci_iswt0;
  output ist_resp_stream_rsci_wen_comp;
  input [106:0] ist_resp_stream_rsci_idat;


  // Interconnect Declarations
  wire ist_resp_stream_rsci_biwt;
  wire ist_resp_stream_rsci_bdwt;
  wire ist_resp_stream_rsci_bcwt;
  wire ist_resp_stream_rsci_irdy;
  wire ist_resp_stream_rsci_ivld_core_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd30),
  .width(32'sd107)) ist_resp_stream_rsci (
      .irdy(ist_resp_stream_rsci_irdy),
      .ivld(ist_resp_stream_rsci_ivld_core_sct),
      .idat(ist_resp_stream_rsci_idat),
      .rdy(ist_resp_stream_rsc_rdy),
      .vld(ist_resp_stream_rsc_vld),
      .dat(ist_resp_stream_rsc_dat)
    );
  ist_core_ist_resp_stream_rsci_ist_resp_stream_wait_ctrl ist_core_ist_resp_stream_rsci_ist_resp_stream_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .ist_resp_stream_rsci_oswt_unreg(ist_resp_stream_rsci_oswt_unreg),
      .ist_resp_stream_rsci_iswt0(ist_resp_stream_rsci_iswt0),
      .ist_resp_stream_rsci_biwt(ist_resp_stream_rsci_biwt),
      .ist_resp_stream_rsci_bdwt(ist_resp_stream_rsci_bdwt),
      .ist_resp_stream_rsci_bcwt(ist_resp_stream_rsci_bcwt),
      .ist_resp_stream_rsci_irdy(ist_resp_stream_rsci_irdy),
      .ist_resp_stream_rsci_ivld_core_sct(ist_resp_stream_rsci_ivld_core_sct)
    );
  ist_core_ist_resp_stream_rsci_ist_resp_stream_wait_dp ist_core_ist_resp_stream_rsci_ist_resp_stream_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ist_resp_stream_rsci_oswt_unreg(ist_resp_stream_rsci_oswt_unreg),
      .ist_resp_stream_rsci_bawt(ist_resp_stream_rsci_bawt),
      .ist_resp_stream_rsci_wen_comp(ist_resp_stream_rsci_wen_comp),
      .ist_resp_stream_rsci_biwt(ist_resp_stream_rsci_biwt),
      .ist_resp_stream_rsci_bdwt(ist_resp_stream_rsci_bdwt),
      .ist_resp_stream_rsci_bcwt(ist_resp_stream_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core_ist_req_stream_rsci
// ------------------------------------------------------------------


module ist_core_ist_req_stream_rsci (
  clk, arst_n, ist_req_stream_rsc_dat, ist_req_stream_rsc_vld, ist_req_stream_rsc_rdy,
      core_wen, ist_req_stream_rsci_oswt_unreg, ist_req_stream_rsci_bawt, ist_req_stream_rsci_iswt0,
      ist_req_stream_rsci_wen_comp, ist_req_stream_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [553:0] ist_req_stream_rsc_dat;
  input ist_req_stream_rsc_vld;
  output ist_req_stream_rsc_rdy;
  input core_wen;
  input ist_req_stream_rsci_oswt_unreg;
  output ist_req_stream_rsci_bawt;
  input ist_req_stream_rsci_iswt0;
  output ist_req_stream_rsci_wen_comp;
  output [553:0] ist_req_stream_rsci_idat_mxwt;


  // Interconnect Declarations
  wire ist_req_stream_rsci_biwt;
  wire ist_req_stream_rsci_bdwt;
  wire ist_req_stream_rsci_bcwt;
  wire ist_req_stream_rsci_irdy_core_sct;
  wire ist_req_stream_rsci_ivld;
  wire [553:0] ist_req_stream_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd29),
  .width(32'sd554)) ist_req_stream_rsci (
      .rdy(ist_req_stream_rsc_rdy),
      .vld(ist_req_stream_rsc_vld),
      .dat(ist_req_stream_rsc_dat),
      .irdy(ist_req_stream_rsci_irdy_core_sct),
      .ivld(ist_req_stream_rsci_ivld),
      .idat(ist_req_stream_rsci_idat)
    );
  ist_core_ist_req_stream_rsci_ist_req_stream_wait_ctrl ist_core_ist_req_stream_rsci_ist_req_stream_wait_ctrl_inst
      (
      .core_wen(core_wen),
      .ist_req_stream_rsci_oswt_unreg(ist_req_stream_rsci_oswt_unreg),
      .ist_req_stream_rsci_iswt0(ist_req_stream_rsci_iswt0),
      .ist_req_stream_rsci_biwt(ist_req_stream_rsci_biwt),
      .ist_req_stream_rsci_bdwt(ist_req_stream_rsci_bdwt),
      .ist_req_stream_rsci_bcwt(ist_req_stream_rsci_bcwt),
      .ist_req_stream_rsci_irdy_core_sct(ist_req_stream_rsci_irdy_core_sct),
      .ist_req_stream_rsci_ivld(ist_req_stream_rsci_ivld)
    );
  ist_core_ist_req_stream_rsci_ist_req_stream_wait_dp ist_core_ist_req_stream_rsci_ist_req_stream_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .ist_req_stream_rsci_oswt_unreg(ist_req_stream_rsci_oswt_unreg),
      .ist_req_stream_rsci_bawt(ist_req_stream_rsci_bawt),
      .ist_req_stream_rsci_wen_comp(ist_req_stream_rsci_wen_comp),
      .ist_req_stream_rsci_idat_mxwt(ist_req_stream_rsci_idat_mxwt),
      .ist_req_stream_rsci_biwt(ist_req_stream_rsci_biwt),
      .ist_req_stream_rsci_bdwt(ist_req_stream_rsci_bdwt),
      .ist_req_stream_rsci_bcwt(ist_req_stream_rsci_bcwt),
      .ist_req_stream_rsci_idat(ist_req_stream_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    init_core
// ------------------------------------------------------------------


module init_core (
  clk, arst_n, init_req_stream_rsc_dat, init_req_stream_rsc_vld, init_req_stream_rsc_rdy,
      trv_req_stream_rsc_dat, trv_req_stream_rsc_vld, trv_req_stream_rsc_rdy
);
  input clk;
  input arst_n;
  input [361:0] init_req_stream_rsc_dat;
  input init_req_stream_rsc_vld;
  output init_req_stream_rsc_rdy;
  output [457:0] trv_req_stream_rsc_dat;
  output trv_req_stream_rsc_vld;
  input trv_req_stream_rsc_rdy;


  // Interconnect Declarations
  wire core_wen;
  wire core_wten;
  wire init_req_stream_rsci_bawt;
  reg init_req_stream_rsci_iswt0;
  wire init_req_stream_rsci_wen_comp;
  wire [361:0] init_req_stream_rsci_idat_mxwt;
  wire trv_req_stream_rsci_bawt;
  wire trv_req_stream_rsci_wen_comp;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt;
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_bawt;
  wire [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_z_mxwt;
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_1_bawt;
  wire [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_1_z_mxwt;
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_2_bawt;
  wire [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_2_z_mxwt;
  reg [63:0] trv_req_stream_rsci_idat_457_394;
  reg [31:0] trv_req_stream_rsci_idat_393_362;
  reg [31:0] trv_req_stream_rsci_idat_361_330;
  reg [31:0] trv_req_stream_rsci_idat_329_298;
  reg [31:0] trv_req_stream_rsci_idat_297_266;
  reg [31:0] trv_req_stream_rsci_idat_265_234;
  reg [31:0] trv_req_stream_rsci_idat_233_202;
  reg [201:0] trv_req_stream_rsci_idat_201_0;
  wire [1:0] fsm_output;
  wire and_11_tmp;
  wire and_9_tmp;
  wire and_7_tmp;
  wire or_dcpl_5;
  wire or_dcpl_6;
  wire or_dcpl_7;
  wire and_dcpl_9;
  wire and_dcpl_10;
  wire and_dcpl_11;
  wire and_dcpl_13;
  reg main_stage_v_3;
  wire or_1_cse_1;
  wire or_2_cse_1;
  wire or_3_cse_1;
  wire or_cse_1;
  reg main_stage_v_4;
  wire and_87_cse;
  reg reg_ccs_lp_piped_fp_recip_23_8_0_cmp_2_iswt1_cse;
  reg reg_ccs_lp_piped_fp_recip_23_8_0_cmp_2_oswt_cse;
  wire init_req_stream_ray_tmax_d_and_2_cse;
  wire init_req_stream_ray_tmax_d_and_3_cse;
  wire and_cse;
  reg reg_trv_req_stream_rsci_iswt0_cse;
  wire and_102_cse;
  wire and_104_cse;
  wire and_103_cse;
  reg main_stage_v_1;
  reg main_stage_v_2;
  reg [31:0] w_x_d_sva_1;
  reg [31:0] w_x_d_sva_2;
  reg [31:0] w_y_d_sva_1;
  reg [31:0] w_y_d_sva_2;
  reg [31:0] w_z_d_sva_1;
  reg [31:0] w_z_d_sva_2;
  reg [63:0] init_req_stream_ray_tmax_d_slc_init_req_stream_crt_265_234_itm_1;
  reg [63:0] init_req_stream_ray_tmax_d_slc_init_req_stream_crt_265_234_itm_2;
  reg [63:0] init_req_stream_ray_tmax_d_slc_init_req_stream_crt_265_234_itm_3;
  reg [63:0] init_req_stream_ray_tmax_d_slc_init_req_stream_crt_265_234_itm_4;
  reg [201:0] init_req_stream_ray_dir_z_d_slc_init_req_stream_crt_201_170_itm_1;
  reg [201:0] init_req_stream_ray_dir_z_d_slc_init_req_stream_crt_201_170_itm_2;
  reg [201:0] init_req_stream_ray_dir_z_d_slc_init_req_stream_crt_201_170_itm_3;
  reg [201:0] init_req_stream_ray_dir_z_d_slc_init_req_stream_crt_201_170_itm_4;
  wire main_stage_v_3_mx0c1;
  wire main_stage_v_4_mx0c1;
  wire main_stage_v_2_mx0c1;
  wire main_stage_v_1_mx0c1;
  wire or_9_cse_1;
  wire or_10_cse_1;
  wire or_11_cse_1;
  wire or_12_cse_1;
  wire or_13_cse_1;
  wire or_14_cse_1;
  wire init_req_stream_ray_tmax_d_and_4_cse;
  wire w_x_d_and_2_cse;

  wire mux_16_nl;
  wire and_114_nl;
  wire or_15_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [457:0] nl_init_core_trv_req_stream_rsci_inst_trv_req_stream_rsci_idat;
  assign nl_init_core_trv_req_stream_rsci_inst_trv_req_stream_rsci_idat = {trv_req_stream_rsci_idat_457_394
      , trv_req_stream_rsci_idat_393_362 , trv_req_stream_rsci_idat_361_330 , trv_req_stream_rsci_idat_329_298
      , trv_req_stream_rsci_idat_297_266 , trv_req_stream_rsci_idat_265_234 , trv_req_stream_rsci_idat_233_202
      , trv_req_stream_rsci_idat_201_0};
  wire [31:0] nl_init_core_ccs_lp_piped_fp_add_23_8_0_cmp_inst_ccs_lp_piped_fp_add_23_8_0_cmp_a_core;
  assign nl_init_core_ccs_lp_piped_fp_add_23_8_0_cmp_inst_ccs_lp_piped_fp_add_23_8_0_cmp_a_core
      = init_req_stream_rsci_idat_mxwt[297:266];
  wire [31:0] nl_init_core_ccs_lp_piped_fp_add_23_8_0_cmp_inst_ccs_lp_piped_fp_add_23_8_0_cmp_b_core;
  assign nl_init_core_ccs_lp_piped_fp_add_23_8_0_cmp_inst_ccs_lp_piped_fp_add_23_8_0_cmp_b_core
      = {(~ (init_req_stream_rsci_idat_mxwt[41])) , (init_req_stream_rsci_idat_mxwt[40:10])};
  wire [31:0] nl_init_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_inst_ccs_lp_piped_fp_add_23_8_0_cmp_1_a_core;
  assign nl_init_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_inst_ccs_lp_piped_fp_add_23_8_0_cmp_1_a_core
      = init_req_stream_rsci_idat_mxwt[361:330];
  wire [31:0] nl_init_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_inst_ccs_lp_piped_fp_add_23_8_0_cmp_1_b_core;
  assign nl_init_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_inst_ccs_lp_piped_fp_add_23_8_0_cmp_1_b_core
      = {(~ (init_req_stream_rsci_idat_mxwt[105])) , (init_req_stream_rsci_idat_mxwt[104:74])};
  wire [31:0] nl_init_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_inst_ccs_lp_piped_fp_add_23_8_0_cmp_2_a_core;
  assign nl_init_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_inst_ccs_lp_piped_fp_add_23_8_0_cmp_2_a_core
      = init_req_stream_rsci_idat_mxwt[329:298];
  wire [31:0] nl_init_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_inst_ccs_lp_piped_fp_add_23_8_0_cmp_2_b_core;
  assign nl_init_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_inst_ccs_lp_piped_fp_add_23_8_0_cmp_2_b_core
      = {(~ (init_req_stream_rsci_idat_mxwt[73])) , (init_req_stream_rsci_idat_mxwt[72:42])};
  wire [31:0] nl_init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_inst_ccs_lp_piped_fp_recip_23_8_0_cmp_a_core;
  assign nl_init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_inst_ccs_lp_piped_fp_recip_23_8_0_cmp_a_core
      = init_req_stream_rsci_idat_mxwt[137:106];
  wire [31:0] nl_init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_1_inst_ccs_lp_piped_fp_recip_23_8_0_cmp_1_a_core;
  assign nl_init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_1_inst_ccs_lp_piped_fp_recip_23_8_0_cmp_1_a_core
      = init_req_stream_rsci_idat_mxwt[201:170];
  wire [31:0] nl_init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_2_inst_ccs_lp_piped_fp_recip_23_8_0_cmp_2_a_core;
  assign nl_init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_2_inst_ccs_lp_piped_fp_recip_23_8_0_cmp_2_a_core
      = init_req_stream_rsci_idat_mxwt[169:138];
  wire  nl_init_core_staller_inst_core_flen_unreg;
  assign nl_init_core_staller_inst_core_flen_unreg = ~((~((~ and_11_tmp) & (fsm_output[1])))
      | and_102_cse | and_103_cse | and_104_cse | (main_stage_v_3 & (~(main_stage_v_4
      & or_dcpl_7)) & or_1_cse_1 & or_2_cse_1 & or_3_cse_1 & or_cse_1 & (fsm_output[1]))
      | (main_stage_v_4 & (~(reg_trv_req_stream_rsci_iswt0_cse & (~ trv_req_stream_rsci_bawt)))
      & or_1_cse_1 & or_2_cse_1 & or_3_cse_1 & or_cse_1 & (fsm_output[1])) | (reg_trv_req_stream_rsci_iswt0_cse
      & or_cse_1 & (fsm_output[1])));
  init_core_init_req_stream_rsci init_core_init_req_stream_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .init_req_stream_rsc_dat(init_req_stream_rsc_dat),
      .init_req_stream_rsc_vld(init_req_stream_rsc_vld),
      .init_req_stream_rsc_rdy(init_req_stream_rsc_rdy),
      .core_wen(core_wen),
      .init_req_stream_rsci_oswt_unreg(and_102_cse),
      .init_req_stream_rsci_bawt(init_req_stream_rsci_bawt),
      .init_req_stream_rsci_iswt0(init_req_stream_rsci_iswt0),
      .init_req_stream_rsci_wen_comp(init_req_stream_rsci_wen_comp),
      .init_req_stream_rsci_idat_mxwt(init_req_stream_rsci_idat_mxwt)
    );
  init_core_trv_req_stream_rsci init_core_trv_req_stream_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .trv_req_stream_rsc_dat(trv_req_stream_rsc_dat),
      .trv_req_stream_rsc_vld(trv_req_stream_rsc_vld),
      .trv_req_stream_rsc_rdy(trv_req_stream_rsc_rdy),
      .core_wen(core_wen),
      .trv_req_stream_rsci_oswt_unreg(and_dcpl_10),
      .trv_req_stream_rsci_bawt(trv_req_stream_rsci_bawt),
      .trv_req_stream_rsci_iswt0(reg_trv_req_stream_rsci_iswt0_cse),
      .trv_req_stream_rsci_wen_comp(trv_req_stream_rsci_wen_comp),
      .trv_req_stream_rsci_idat(nl_init_core_trv_req_stream_rsci_inst_trv_req_stream_rsci_idat[457:0])
    );
  init_core_ccs_lp_piped_fp_mult_23_8_0_cmp init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_oswt_unreg(and_dcpl_9),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1(reg_ccs_lp_piped_fp_recip_23_8_0_cmp_2_oswt_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_a_core(ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_b_core(ccs_lp_piped_fp_recip_23_8_0_cmp_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1_pff(and_104_cse)
    );
  init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1 init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_oswt_unreg(and_dcpl_9),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1(reg_ccs_lp_piped_fp_recip_23_8_0_cmp_2_oswt_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_a_core(ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_b_core(ccs_lp_piped_fp_recip_23_8_0_cmp_1_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1_pff(and_104_cse)
    );
  init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2 init_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_oswt_unreg(and_dcpl_9),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1(reg_ccs_lp_piped_fp_recip_23_8_0_cmp_2_oswt_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_a_core(ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_b_core(ccs_lp_piped_fp_recip_23_8_0_cmp_2_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1_pff(and_104_cse)
    );
  init_core_ccs_lp_piped_fp_add_23_8_0_cmp init_core_ccs_lp_piped_fp_add_23_8_0_cmp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_oswt_unreg(and_104_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_iswt1(reg_ccs_lp_piped_fp_recip_23_8_0_cmp_2_iswt1_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_a_core(nl_init_core_ccs_lp_piped_fp_add_23_8_0_cmp_inst_ccs_lp_piped_fp_add_23_8_0_cmp_a_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_b_core(nl_init_core_ccs_lp_piped_fp_add_23_8_0_cmp_inst_ccs_lp_piped_fp_add_23_8_0_cmp_b_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_iswt1_pff(and_102_cse)
    );
  init_core_ccs_lp_piped_fp_add_23_8_0_cmp_1 init_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_oswt_unreg(and_104_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1(reg_ccs_lp_piped_fp_recip_23_8_0_cmp_2_iswt1_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_a_core(nl_init_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_inst_ccs_lp_piped_fp_add_23_8_0_cmp_1_a_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_b_core(nl_init_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_inst_ccs_lp_piped_fp_add_23_8_0_cmp_1_b_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1_pff(and_102_cse)
    );
  init_core_ccs_lp_piped_fp_add_23_8_0_cmp_2 init_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_oswt_unreg(and_104_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1(reg_ccs_lp_piped_fp_recip_23_8_0_cmp_2_iswt1_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_a_core(nl_init_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_inst_ccs_lp_piped_fp_add_23_8_0_cmp_2_a_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_b_core(nl_init_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_inst_ccs_lp_piped_fp_add_23_8_0_cmp_2_b_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1_pff(and_102_cse)
    );
  init_core_ccs_lp_piped_fp_recip_23_8_0_cmp init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_oswt_unreg(and_104_cse),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_bawt(ccs_lp_piped_fp_recip_23_8_0_cmp_bawt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1(reg_ccs_lp_piped_fp_recip_23_8_0_cmp_2_iswt1_cse),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_a_core(nl_init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_inst_ccs_lp_piped_fp_recip_23_8_0_cmp_a_core[31:0]),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_z_mxwt(ccs_lp_piped_fp_recip_23_8_0_cmp_z_mxwt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1_pff(and_102_cse)
    );
  init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_1 init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_1_oswt_unreg(and_104_cse),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_1_bawt(ccs_lp_piped_fp_recip_23_8_0_cmp_1_bawt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_1_iswt1(reg_ccs_lp_piped_fp_recip_23_8_0_cmp_2_iswt1_cse),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_1_a_core(nl_init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_1_inst_ccs_lp_piped_fp_recip_23_8_0_cmp_1_a_core[31:0]),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_1_z_mxwt(ccs_lp_piped_fp_recip_23_8_0_cmp_1_z_mxwt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_1_iswt1_pff(and_102_cse)
    );
  init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_2 init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_2_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_2_oswt_unreg(and_104_cse),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_2_bawt(ccs_lp_piped_fp_recip_23_8_0_cmp_2_bawt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_2_iswt1(reg_ccs_lp_piped_fp_recip_23_8_0_cmp_2_iswt1_cse),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_2_a_core(nl_init_core_ccs_lp_piped_fp_recip_23_8_0_cmp_2_inst_ccs_lp_piped_fp_recip_23_8_0_cmp_2_a_core[31:0]),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_2_z_mxwt(ccs_lp_piped_fp_recip_23_8_0_cmp_2_z_mxwt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_2_iswt1_pff(and_102_cse)
    );
  init_core_staller init_core_staller_inst (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .init_req_stream_rsci_wen_comp(init_req_stream_rsci_wen_comp),
      .trv_req_stream_rsci_wen_comp(trv_req_stream_rsci_wen_comp),
      .core_flen_unreg(nl_init_core_staller_inst_core_flen_unreg)
    );
  init_core_core_fsm init_core_core_fsm_inst (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign and_87_cse = core_wen & (~ or_dcpl_7);
  assign and_102_cse = and_11_tmp & (fsm_output[1]);
  assign and_104_cse = and_7_tmp & (fsm_output[1]);
  assign and_103_cse = and_9_tmp & (fsm_output[1]);
  assign and_114_nl = main_stage_v_4 & (~(or_cse_1 & ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt
      & ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt & ccs_lp_piped_fp_mult_23_8_0_cmp_bawt));
  assign or_15_nl = main_stage_v_4 | (~ reg_trv_req_stream_rsci_iswt0_cse) | trv_req_stream_rsci_bawt;
  assign mux_16_nl = MUX_s_1_2_2(and_114_nl, or_15_nl, main_stage_v_3);
  assign init_req_stream_ray_tmax_d_and_4_cse = core_wen & (~((or_dcpl_6 & main_stage_v_4)
      | and_cse)) & mux_16_nl;
  assign w_x_d_and_2_cse = core_wen & and_7_tmp;
  assign init_req_stream_ray_tmax_d_and_2_cse = core_wen & (~((~ and_9_tmp) | (fsm_output[0])));
  assign init_req_stream_ray_tmax_d_and_3_cse = core_wen & (~((~ and_11_tmp) | (fsm_output[0])));
  assign and_11_tmp = init_req_stream_rsci_bawt & or_9_cse_1 & or_10_cse_1 & or_11_cse_1
      & or_12_cse_1 & or_13_cse_1 & or_14_cse_1 & or_1_cse_1 & or_2_cse_1 & or_3_cse_1
      & or_cse_1;
  assign and_9_tmp = main_stage_v_1 & or_9_cse_1 & or_10_cse_1 & or_11_cse_1 & or_12_cse_1
      & or_13_cse_1 & or_14_cse_1 & or_1_cse_1 & or_2_cse_1 & or_3_cse_1 & or_cse_1;
  assign and_7_tmp = main_stage_v_2 & or_9_cse_1 & or_10_cse_1 & or_11_cse_1 & or_12_cse_1
      & or_13_cse_1 & or_14_cse_1 & or_1_cse_1 & or_2_cse_1 & or_3_cse_1 & or_cse_1;
  assign or_9_cse_1 = ccs_lp_piped_fp_recip_23_8_0_cmp_bawt | (~ main_stage_v_2);
  assign or_10_cse_1 = ccs_lp_piped_fp_recip_23_8_0_cmp_2_bawt | (~ main_stage_v_2);
  assign or_11_cse_1 = ccs_lp_piped_fp_recip_23_8_0_cmp_1_bawt | (~ main_stage_v_2);
  assign or_12_cse_1 = ccs_lp_piped_fp_add_23_8_0_cmp_bawt | (~ main_stage_v_2);
  assign or_13_cse_1 = ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt | (~ main_stage_v_2);
  assign or_14_cse_1 = ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt | (~ main_stage_v_2);
  assign or_1_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_bawt | (~ main_stage_v_4);
  assign or_2_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt | (~ main_stage_v_4);
  assign or_3_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt | (~ main_stage_v_4);
  assign or_cse_1 = trv_req_stream_rsci_bawt | (~ reg_trv_req_stream_rsci_iswt0_cse);
  assign and_cse = (~ trv_req_stream_rsci_bawt) & reg_trv_req_stream_rsci_iswt0_cse;
  assign or_dcpl_5 = ~(ccs_lp_piped_fp_mult_23_8_0_cmp_bawt & ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt);
  assign or_dcpl_6 = or_dcpl_5 | (~ ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt);
  assign or_dcpl_7 = or_dcpl_6 | and_cse | (~ main_stage_v_4);
  assign and_dcpl_9 = or_cse_1 & ccs_lp_piped_fp_mult_23_8_0_cmp_bawt & ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt
      & ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt & main_stage_v_4;
  assign and_dcpl_10 = trv_req_stream_rsci_bawt & reg_trv_req_stream_rsci_iswt0_cse;
  assign and_dcpl_11 = (or_dcpl_5 | (~(ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt & main_stage_v_4)))
      & and_dcpl_10;
  assign and_dcpl_13 = (~((~(ccs_lp_piped_fp_mult_23_8_0_cmp_bawt & ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt
      & ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt)) & main_stage_v_4)) & or_cse_1;
  assign main_stage_v_3_mx0c1 = and_dcpl_13 & main_stage_v_3 & (~ and_7_tmp);
  assign main_stage_v_4_mx0c1 = ccs_lp_piped_fp_mult_23_8_0_cmp_bawt & ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt
      & or_cse_1 & ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt & main_stage_v_4 & (~ main_stage_v_3);
  assign main_stage_v_2_mx0c1 = and_7_tmp & (~ and_9_tmp) & (fsm_output[1]);
  assign main_stage_v_1_mx0c1 = and_9_tmp & (~ and_11_tmp) & (fsm_output[1]);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      init_req_stream_rsci_iswt0 <= 1'b0;
    end
    else if ( core_wen & (and_11_tmp | (fsm_output[0])) ) begin
      init_req_stream_rsci_iswt0 <= 1'b1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      trv_req_stream_rsci_idat_201_0 <= 202'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      trv_req_stream_rsci_idat_233_202 <= 32'b00000000000000000000000000000000;
      trv_req_stream_rsci_idat_265_234 <= 32'b00000000000000000000000000000000;
      trv_req_stream_rsci_idat_297_266 <= 32'b00000000000000000000000000000000;
      trv_req_stream_rsci_idat_329_298 <= 32'b00000000000000000000000000000000;
      trv_req_stream_rsci_idat_361_330 <= 32'b00000000000000000000000000000000;
      trv_req_stream_rsci_idat_393_362 <= 32'b00000000000000000000000000000000;
      trv_req_stream_rsci_idat_457_394 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_87_cse ) begin
      trv_req_stream_rsci_idat_201_0 <= init_req_stream_ray_dir_z_d_slc_init_req_stream_crt_201_170_itm_4;
      trv_req_stream_rsci_idat_233_202 <= w_x_d_sva_2;
      trv_req_stream_rsci_idat_265_234 <= w_y_d_sva_2;
      trv_req_stream_rsci_idat_297_266 <= w_z_d_sva_2;
      trv_req_stream_rsci_idat_329_298 <= ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt;
      trv_req_stream_rsci_idat_361_330 <= ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt;
      trv_req_stream_rsci_idat_393_362 <= ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt;
      trv_req_stream_rsci_idat_457_394 <= init_req_stream_ray_tmax_d_slc_init_req_stream_crt_265_234_itm_4;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_ccs_lp_piped_fp_recip_23_8_0_cmp_2_iswt1_cse <= 1'b0;
      reg_ccs_lp_piped_fp_recip_23_8_0_cmp_2_oswt_cse <= 1'b0;
    end
    else if ( core_wen ) begin
      reg_ccs_lp_piped_fp_recip_23_8_0_cmp_2_iswt1_cse <= and_102_cse;
      reg_ccs_lp_piped_fp_recip_23_8_0_cmp_2_oswt_cse <= and_104_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_trv_req_stream_rsci_iswt0_cse <= 1'b0;
    end
    else if ( core_wen & (and_dcpl_9 | and_dcpl_11) ) begin
      reg_trv_req_stream_rsci_iswt0_cse <= ~ and_dcpl_11;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_3 <= 1'b0;
    end
    else if ( core_wen & (and_104_cse | main_stage_v_3_mx0c1) ) begin
      main_stage_v_3 <= ~ main_stage_v_3_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_4 <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_13 & main_stage_v_3) | main_stage_v_4_mx0c1)
        ) begin
      main_stage_v_4 <= ~ main_stage_v_4_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      init_req_stream_ray_tmax_d_slc_init_req_stream_crt_265_234_itm_4 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      init_req_stream_ray_dir_z_d_slc_init_req_stream_crt_201_170_itm_4 <= 202'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      w_x_d_sva_2 <= 32'b00000000000000000000000000000000;
      w_y_d_sva_2 <= 32'b00000000000000000000000000000000;
      w_z_d_sva_2 <= 32'b00000000000000000000000000000000;
    end
    else if ( init_req_stream_ray_tmax_d_and_4_cse ) begin
      init_req_stream_ray_tmax_d_slc_init_req_stream_crt_265_234_itm_4 <= init_req_stream_ray_tmax_d_slc_init_req_stream_crt_265_234_itm_3;
      init_req_stream_ray_dir_z_d_slc_init_req_stream_crt_201_170_itm_4 <= init_req_stream_ray_dir_z_d_slc_init_req_stream_crt_201_170_itm_3;
      w_x_d_sva_2 <= w_x_d_sva_1;
      w_y_d_sva_2 <= w_y_d_sva_1;
      w_z_d_sva_2 <= w_z_d_sva_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_2 <= 1'b0;
    end
    else if ( core_wen & (and_103_cse | main_stage_v_2_mx0c1) ) begin
      main_stage_v_2 <= ~ main_stage_v_2_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_1 <= 1'b0;
    end
    else if ( core_wen & (and_102_cse | main_stage_v_1_mx0c1) ) begin
      main_stage_v_1 <= ~ main_stage_v_1_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      w_x_d_sva_1 <= 32'b00000000000000000000000000000000;
      w_y_d_sva_1 <= 32'b00000000000000000000000000000000;
      w_z_d_sva_1 <= 32'b00000000000000000000000000000000;
      init_req_stream_ray_tmax_d_slc_init_req_stream_crt_265_234_itm_3 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      init_req_stream_ray_dir_z_d_slc_init_req_stream_crt_201_170_itm_3 <= 202'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( w_x_d_and_2_cse ) begin
      w_x_d_sva_1 <= ccs_lp_piped_fp_recip_23_8_0_cmp_z_mxwt;
      w_y_d_sva_1 <= ccs_lp_piped_fp_recip_23_8_0_cmp_2_z_mxwt;
      w_z_d_sva_1 <= ccs_lp_piped_fp_recip_23_8_0_cmp_1_z_mxwt;
      init_req_stream_ray_tmax_d_slc_init_req_stream_crt_265_234_itm_3 <= init_req_stream_ray_tmax_d_slc_init_req_stream_crt_265_234_itm_2;
      init_req_stream_ray_dir_z_d_slc_init_req_stream_crt_201_170_itm_3 <= init_req_stream_ray_dir_z_d_slc_init_req_stream_crt_201_170_itm_2;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      init_req_stream_ray_tmax_d_slc_init_req_stream_crt_265_234_itm_2 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      init_req_stream_ray_dir_z_d_slc_init_req_stream_crt_201_170_itm_2 <= 202'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( init_req_stream_ray_tmax_d_and_2_cse ) begin
      init_req_stream_ray_tmax_d_slc_init_req_stream_crt_265_234_itm_2 <= init_req_stream_ray_tmax_d_slc_init_req_stream_crt_265_234_itm_1;
      init_req_stream_ray_dir_z_d_slc_init_req_stream_crt_201_170_itm_2 <= init_req_stream_ray_dir_z_d_slc_init_req_stream_crt_201_170_itm_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      init_req_stream_ray_tmax_d_slc_init_req_stream_crt_265_234_itm_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      init_req_stream_ray_dir_z_d_slc_init_req_stream_crt_201_170_itm_1 <= 202'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( init_req_stream_ray_tmax_d_and_3_cse ) begin
      init_req_stream_ray_tmax_d_slc_init_req_stream_crt_265_234_itm_1 <= init_req_stream_rsci_idat_mxwt[265:202];
      init_req_stream_ray_dir_z_d_slc_init_req_stream_crt_201_170_itm_1 <= init_req_stream_rsci_idat_mxwt[201:0];
    end
  end

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox_core
// ------------------------------------------------------------------


module bbox_core (
  clk, arst_n, bbox_req_stream_rsc_dat, bbox_req_stream_rsc_vld, bbox_req_stream_rsc_rdy,
      bbox_resp_stream_rsc_dat, bbox_resp_stream_rsc_vld, bbox_resp_stream_rsc_rdy
);
  input clk;
  input arst_n;
  input [385:0] bbox_req_stream_rsc_dat;
  input bbox_req_stream_rsc_vld;
  output bbox_req_stream_rsc_rdy;
  output [204:0] bbox_resp_stream_rsc_dat;
  output bbox_resp_stream_rsc_vld;
  input bbox_resp_stream_rsc_rdy;


  // Interconnect Declarations
  wire core_wen;
  wire core_wten;
  wire bbox_req_stream_rsci_bawt;
  reg bbox_req_stream_rsci_iswt0;
  wire bbox_req_stream_rsci_wen_comp;
  wire [385:0] bbox_req_stream_rsci_idat_mxwt;
  wire bbox_resp_stream_rsci_bawt;
  wire bbox_resp_stream_rsci_wen_comp;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_3_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_3_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_4_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_4_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_5_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_5_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_6_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_6_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_7_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_7_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_8_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_8_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_9_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_9_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_10_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_10_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_11_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_11_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_3_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_5_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_6_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_7_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_8_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_9_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_10_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_11_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_12_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_13_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_14_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_15_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_16_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_17_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_18_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_19_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_20_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_21_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_22_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_23_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_mxwt;
  reg bbox_resp_stream_rsci_idat_204;
  reg bbox_resp_stream_rsci_idat_203;
  reg bbox_resp_stream_rsci_idat_202;
  reg [31:0] bbox_resp_stream_rsci_idat_201_170;
  reg [31:0] bbox_resp_stream_rsci_idat_169_138;
  reg [31:0] bbox_resp_stream_rsci_idat_137_106;
  reg [31:0] bbox_resp_stream_rsci_idat_105_74;
  reg [31:0] bbox_resp_stream_rsci_idat_73_42;
  reg [31:0] bbox_resp_stream_rsci_idat_41_10;
  reg [9:0] bbox_resp_stream_rsci_idat_9_0;
  wire [1:0] fsm_output;
  wire and_17_tmp;
  wire and_15_tmp;
  wire and_13_tmp;
  wire and_11_tmp;
  wire and_9_tmp;
  wire and_7_tmp;
  wire and_5_tmp;
  wire and_dcpl_6;
  wire and_dcpl_7;
  wire and_dcpl_12;
  wire and_dcpl_14;
  wire and_dcpl_16;
  wire [7:0] bbox_ns_ldexpf_a_11_lpi_1_dfm_mx0;
  wire [7:0] bbox_ns_ldexpf_a_10_lpi_1_dfm_mx0;
  wire [7:0] bbox_ns_ldexpf_a_9_lpi_1_dfm_mx0;
  wire [7:0] bbox_ns_ldexpf_a_8_lpi_1_dfm_mx0;
  wire [7:0] bbox_ns_ldexpf_a_7_lpi_1_dfm_mx0;
  wire [7:0] bbox_ns_ldexpf_a_6_lpi_1_dfm_mx0;
  wire [7:0] bbox_ns_ldexpf_a_5_lpi_1_dfm_mx0;
  wire [7:0] bbox_ns_ldexpf_a_4_lpi_1_dfm_mx0;
  wire [7:0] bbox_ns_ldexpf_a_3_lpi_1_dfm_mx0;
  wire [7:0] bbox_ns_ldexpf_a_2_lpi_1_dfm_mx0;
  wire [7:0] bbox_ns_ldexpf_a_1_lpi_1_dfm_mx0;
  wire [7:0] bbox_ns_ldexpf_a_lpi_1_dfm_mx0;
  reg main_stage_v_7;
  wire or_cse_1;
  reg bbox_req_stream_crt_sva_6_41;
  reg bbox_req_stream_crt_sva_6_73;
  reg bbox_req_stream_crt_sva_6_105;
  wire and_169_cse;
  reg reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1_cse;
  reg reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_cse;
  reg reg_ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1_cse;
  wire and_192_cse;
  wire and_199_cse;
  wire and_187_cse;
  wire and_197_cse;
  reg reg_bbox_resp_stream_rsci_iswt0_cse;
  wire and_213_cse;
  wire and_215_cse;
  wire and_211_cse;
  wire and_217_cse;
  wire and_216_cse;
  wire and_214_cse;
  wire and_212_cse;
  wire [7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_x_u_sva_1;
  wire [7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_11_x_u_sva_1;
  wire [7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_10_x_u_sva_1;
  wire [7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_9_x_u_sva_1;
  wire [7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_8_x_u_sva_1;
  wire [7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_7_x_u_sva_1;
  wire [7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_6_x_u_sva_1;
  wire [7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_5_x_u_sva_1;
  wire [7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_4_x_u_sva_1;
  wire [7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_3_x_u_sva_1;
  wire [7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_2_x_u_sva_1;
  wire [7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_1_x_u_sva_1;
  reg [160:0] bbox_req_stream_crt_sva_4_265_105;
  reg [265:0] bbox_req_stream_crt_sva_2_265_0;
  reg [63:0] bbox_req_stream_crt_sva_6_265_202;
  wire [7:0] status0_out;
  wire [7:0] status1_out;
  wire [7:0] status0_out_1;
  wire [7:0] status1_out_1;
  wire [7:0] status0_out_2;
  wire [7:0] status1_out_2;
  wire [7:0] status0_out_3;
  wire [7:0] status1_out_3;
  wire [7:0] status0_out_4;
  wire [7:0] status1_out_4;
  wire [7:0] status0_out_5;
  wire [7:0] status1_out_5;
  wire [7:0] status0_out_6;
  wire [7:0] status1_out_6;
  wire [7:0] status0_out_7;
  wire [7:0] status1_out_7;
  wire [7:0] status0_out_8;
  wire [7:0] status1_out_8;
  wire [7:0] status0_out_9;
  wire [7:0] status1_out_9;
  wire [7:0] status0_out_10;
  wire [7:0] status1_out_10;
  wire [7:0] status0_out_11;
  wire [7:0] status1_out_11;
  wire [7:0] status0_out_12;
  wire [7:0] status1_out_12;
  wire [7:0] status0_out_13;
  wire [7:0] status1_out_13;
  wire [7:0] status0_out_14;
  wire [7:0] status1_out_14;
  reg main_stage_v_1;
  reg main_stage_v_2;
  reg main_stage_v_3;
  reg main_stage_v_4;
  reg main_stage_v_5;
  reg main_stage_v_6;
  reg [31:0] bbox_ns_fmax_return_d_2_lpi_1_dfm_1;
  reg [31:0] bbox_ns_fmax_return_d_5_lpi_1_dfm_1;
  reg [31:0] return_ac_std_float_23_mux_itm_1;
  reg [31:0] return_ac_std_float_47_mux_itm_1;
  reg [31:0] const_z_min_ac_std_float_1_mux_3_itm_1;
  reg [31:0] const_z_min_ac_std_float_1_mux_2_itm_1;
  reg [31:0] const_x_min_ac_std_float_1_mux_1_itm_1;
  reg [31:0] const_z_min_ac_std_float_1_mux_1_itm_1;
  reg [31:0] const_z_min_ac_std_float_1_mux_itm_1;
  reg [31:0] const_x_min_ac_std_float_1_mux_itm_1;
  reg [9:0] bbox_req_stream_rid_slc_bbox_req_stream_crt_9_0_itm_1;
  reg [265:0] bbox_req_stream_crt_sva_1_265_0;
  reg [160:0] bbox_req_stream_crt_sva_3_265_105;
  reg bbox_req_stream_crt_sva_3_73;
  reg bbox_req_stream_crt_sva_3_41;
  reg [9:0] bbox_req_stream_crt_sva_3_9_0;
  reg bbox_req_stream_crt_sva_4_73;
  reg bbox_req_stream_crt_sva_4_41;
  reg [9:0] bbox_req_stream_crt_sva_4_9_0;
  reg [63:0] bbox_req_stream_crt_sva_5_265_202;
  reg bbox_req_stream_crt_sva_5_105;
  reg bbox_req_stream_crt_sva_5_73;
  reg bbox_req_stream_crt_sva_5_41;
  reg [9:0] bbox_req_stream_crt_sva_5_9_0;
  reg [9:0] bbox_req_stream_crt_sva_6_9_0;
  wire main_stage_v_7_mx0c1;
  wire main_stage_v_6_mx0c1;
  wire main_stage_v_5_mx0c1;
  wire main_stage_v_4_mx0c1;
  wire main_stage_v_3_mx0c1;
  wire main_stage_v_2_mx0c1;
  wire main_stage_v_1_mx0c1;
  wire or_78_cse_1;
  wire or_79_cse_1;
  wire or_80_cse_1;
  wire or_81_cse_1;
  wire or_82_cse_1;
  wire or_83_cse_1;
  wire or_84_cse_1;
  wire or_85_cse_1;
  wire or_86_cse_1;
  wire or_87_cse_1;
  wire or_88_cse_1;
  wire or_89_cse_1;
  wire or_28_cse_1;
  wire or_29_cse_1;
  wire or_30_cse_1;
  wire or_31_cse_1;
  wire or_32_cse_1;
  wire or_33_cse_1;
  wire or_34_cse_1;
  wire or_35_cse_1;
  wire or_36_cse_1;
  wire or_37_cse_1;
  wire or_38_cse_1;
  wire or_39_cse_1;
  wire or_2_cse_1;
  wire or_3_cse_1;
  wire or_4_cse_1;
  wire or_5_cse_1;
  wire or_6_cse_1;
  wire or_7_cse_1;
  wire or_8_cse_1;
  wire or_9_cse_1;
  wire or_10_cse_1;
  wire or_11_cse_1;
  wire or_12_cse_1;
  wire or_13_cse_1;
  wire [31:0] bbox_ns_fmin_return_d_4_lpi_1_dfm_mx0;
  wire [31:0] bbox_ns_fmin_return_d_3_lpi_1_dfm_mx0;
  wire [31:0] bbox_ns_fmax_return_d_3_lpi_1_dfm_mx0;
  wire [31:0] bbox_ns_fmax_return_d_4_lpi_1_dfm_mx0;
  wire [31:0] bbox_ns_fmin_return_d_1_lpi_1_dfm_mx0;
  wire [31:0] bbox_ns_fmin_return_d_lpi_1_dfm_mx0;
  wire [31:0] bbox_ns_fmax_return_d_lpi_1_dfm_mx0;
  wire [31:0] bbox_ns_fmax_return_d_1_lpi_1_dfm_mx0;
  wire ccs_fp_cmp_23_8_0_14_out_6;
  wire ccs_fp_cmp_23_8_0_14_out_7;
  wire ccs_fp_cmp_23_8_0_14_out_8;
  wire ccs_fp_cmp_23_8_0_14_out_9;
  wire [31:0] ccs_fp_cmp_23_8_0_14_out_10;
  wire [31:0] ccs_fp_cmp_23_8_0_14_out_11;
  wire ccs_fp_cmp_23_8_0_13_out_6;
  wire ccs_fp_cmp_23_8_0_13_out_7;
  wire ccs_fp_cmp_23_8_0_13_out_8;
  wire ccs_fp_cmp_23_8_0_13_out_9;
  wire [31:0] ccs_fp_cmp_23_8_0_13_out_10;
  wire [31:0] ccs_fp_cmp_23_8_0_13_out_11;
  wire ccs_fp_cmp_23_8_0_6_out_6;
  wire ccs_fp_cmp_23_8_0_6_out_7;
  wire ccs_fp_cmp_23_8_0_6_out_8;
  wire ccs_fp_cmp_23_8_0_6_out_9;
  wire [31:0] ccs_fp_cmp_23_8_0_6_out_10;
  wire [31:0] ccs_fp_cmp_23_8_0_6_out_11;
  wire [3:0] leading_sign_8_0_1_0_11_out_3;
  wire [3:0] leading_sign_8_0_1_0_10_out_3;
  wire [3:0] leading_sign_8_0_1_0_9_out_3;
  wire [3:0] leading_sign_8_0_1_0_8_out_3;
  wire [3:0] leading_sign_8_0_1_0_7_out_3;
  wire [3:0] leading_sign_8_0_1_0_6_out_3;
  wire [3:0] leading_sign_8_0_1_0_5_out_3;
  wire [3:0] leading_sign_8_0_1_0_4_out_3;
  wire [3:0] leading_sign_8_0_1_0_3_out_3;
  wire [3:0] leading_sign_8_0_1_0_2_out_3;
  wire [3:0] leading_sign_8_0_1_0_1_out_3;
  wire [3:0] leading_sign_8_0_1_0_out_3;
  wire ccs_fp_cmp_23_8_0_12_out_6;
  wire ccs_fp_cmp_23_8_0_12_out_7;
  wire ccs_fp_cmp_23_8_0_12_out_8;
  wire ccs_fp_cmp_23_8_0_12_out_9;
  wire [31:0] ccs_fp_cmp_23_8_0_12_out_10;
  wire [31:0] ccs_fp_cmp_23_8_0_12_out_11;
  wire ccs_fp_cmp_23_8_0_11_out_6;
  wire ccs_fp_cmp_23_8_0_11_out_7;
  wire ccs_fp_cmp_23_8_0_11_out_8;
  wire ccs_fp_cmp_23_8_0_11_out_9;
  wire [31:0] ccs_fp_cmp_23_8_0_11_out_10;
  wire [31:0] ccs_fp_cmp_23_8_0_11_out_11;
  wire ccs_fp_cmp_23_8_0_10_out_6;
  wire ccs_fp_cmp_23_8_0_10_out_7;
  wire ccs_fp_cmp_23_8_0_10_out_8;
  wire ccs_fp_cmp_23_8_0_10_out_9;
  wire [31:0] ccs_fp_cmp_23_8_0_10_out_10;
  wire [31:0] ccs_fp_cmp_23_8_0_10_out_11;
  wire ccs_fp_cmp_23_8_0_9_out_6;
  wire ccs_fp_cmp_23_8_0_9_out_7;
  wire ccs_fp_cmp_23_8_0_9_out_8;
  wire ccs_fp_cmp_23_8_0_9_out_9;
  wire [31:0] ccs_fp_cmp_23_8_0_9_out_10;
  wire [31:0] ccs_fp_cmp_23_8_0_9_out_11;
  wire ccs_fp_cmp_23_8_0_8_out_6;
  wire ccs_fp_cmp_23_8_0_8_out_7;
  wire ccs_fp_cmp_23_8_0_8_out_8;
  wire ccs_fp_cmp_23_8_0_8_out_9;
  wire [31:0] ccs_fp_cmp_23_8_0_8_out_10;
  wire [31:0] ccs_fp_cmp_23_8_0_8_out_11;
  wire ccs_fp_cmp_23_8_0_7_out_6;
  wire ccs_fp_cmp_23_8_0_7_out_7;
  wire ccs_fp_cmp_23_8_0_7_out_8;
  wire ccs_fp_cmp_23_8_0_7_out_9;
  wire [31:0] ccs_fp_cmp_23_8_0_7_out_10;
  wire [31:0] ccs_fp_cmp_23_8_0_7_out_11;
  wire ccs_fp_cmp_23_8_0_5_out_6;
  wire ccs_fp_cmp_23_8_0_5_out_7;
  wire ccs_fp_cmp_23_8_0_5_out_8;
  wire ccs_fp_cmp_23_8_0_5_out_9;
  wire [31:0] ccs_fp_cmp_23_8_0_5_out_10;
  wire [31:0] ccs_fp_cmp_23_8_0_5_out_11;
  wire ccs_fp_cmp_23_8_0_4_out_6;
  wire ccs_fp_cmp_23_8_0_4_out_7;
  wire ccs_fp_cmp_23_8_0_4_out_8;
  wire ccs_fp_cmp_23_8_0_4_out_9;
  wire [31:0] ccs_fp_cmp_23_8_0_4_out_10;
  wire [31:0] ccs_fp_cmp_23_8_0_4_out_11;
  wire ccs_fp_cmp_23_8_0_3_out_6;
  wire ccs_fp_cmp_23_8_0_3_out_7;
  wire ccs_fp_cmp_23_8_0_3_out_8;
  wire ccs_fp_cmp_23_8_0_3_out_9;
  wire [31:0] ccs_fp_cmp_23_8_0_3_out_10;
  wire [31:0] ccs_fp_cmp_23_8_0_3_out_11;
  wire ccs_fp_cmp_23_8_0_2_out_6;
  wire ccs_fp_cmp_23_8_0_2_out_7;
  wire ccs_fp_cmp_23_8_0_2_out_8;
  wire ccs_fp_cmp_23_8_0_2_out_9;
  wire [31:0] ccs_fp_cmp_23_8_0_2_out_10;
  wire [31:0] ccs_fp_cmp_23_8_0_2_out_11;
  wire ccs_fp_cmp_23_8_0_1_out_6;
  wire ccs_fp_cmp_23_8_0_1_out_7;
  wire ccs_fp_cmp_23_8_0_1_out_8;
  wire ccs_fp_cmp_23_8_0_1_out_9;
  wire [31:0] ccs_fp_cmp_23_8_0_1_out_10;
  wire [31:0] ccs_fp_cmp_23_8_0_1_out_11;
  wire ccs_fp_cmp_23_8_0_out_6;
  wire ccs_fp_cmp_23_8_0_out_7;
  wire ccs_fp_cmp_23_8_0_out_8;
  wire ccs_fp_cmp_23_8_0_out_9;
  wire [31:0] ccs_fp_cmp_23_8_0_out_10;
  wire [31:0] ccs_fp_cmp_23_8_0_out_11;
  wire bbox_req_stream_rid_and_1_cse;

  wire and_35_nl;
  wire and_37_nl;
  wire and_39_nl;
  wire and_41_nl;
  wire FP_LEQ_32_8_11_nor_nl;
  wire FP_LEQ_32_8_10_nor_nl;
  wire FP_LEQ_32_8_7_nor_nl;
  wire FP_LEQ_32_8_8_nor_nl;
  wire FP_LEQ_32_8_4_nor_nl;
  wire FP_LEQ_32_8_3_nor_nl;
  wire FP_LEQ_32_8_nor_nl;
  wire FP_LEQ_32_8_1_nor_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_ccs_fp_cmp_23_8_0_11_rg_b;
  assign nl_ccs_fp_cmp_23_8_0_11_rg_b = bbox_req_stream_crt_sva_6_265_202[63:32];
  wire [31:0] nl_ccs_fp_cmp_23_8_0_8_rg_b;
  assign nl_ccs_fp_cmp_23_8_0_8_rg_b = bbox_req_stream_crt_sva_6_265_202[31:0];
  wire [31:0] nl_ccs_fp_cmp_23_8_0_4_rg_b;
  assign nl_ccs_fp_cmp_23_8_0_4_rg_b = bbox_req_stream_crt_sva_6_265_202[63:32];
  wire [31:0] nl_ccs_fp_cmp_23_8_0_1_rg_b;
  assign nl_ccs_fp_cmp_23_8_0_1_rg_b = bbox_req_stream_crt_sva_6_265_202[31:0];
  wire [204:0] nl_bbox_core_bbox_resp_stream_rsci_inst_bbox_resp_stream_rsci_idat;
  assign nl_bbox_core_bbox_resp_stream_rsci_inst_bbox_resp_stream_rsci_idat = {bbox_resp_stream_rsci_idat_204
      , bbox_resp_stream_rsci_idat_203 , bbox_resp_stream_rsci_idat_202 , bbox_resp_stream_rsci_idat_201_170
      , bbox_resp_stream_rsci_idat_169_138 , bbox_resp_stream_rsci_idat_137_106 ,
      bbox_resp_stream_rsci_idat_105_74 , bbox_resp_stream_rsci_idat_73_42 , bbox_resp_stream_rsci_idat_41_10
      , bbox_resp_stream_rsci_idat_9_0};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_inst_ccs_lp_piped_fp_add_23_8_0_cmp_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_inst_ccs_lp_piped_fp_add_23_8_0_cmp_b_core
      = bbox_req_stream_crt_sva_4_265_105[32:1];
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_inst_ccs_lp_piped_fp_add_23_8_0_cmp_1_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_inst_ccs_lp_piped_fp_add_23_8_0_cmp_1_b_core
      = bbox_req_stream_crt_sva_4_265_105[96:65];
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_inst_ccs_lp_piped_fp_add_23_8_0_cmp_2_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_inst_ccs_lp_piped_fp_add_23_8_0_cmp_2_b_core
      = bbox_req_stream_crt_sva_4_265_105[64:33];
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_3_inst_ccs_lp_piped_fp_add_23_8_0_cmp_3_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_3_inst_ccs_lp_piped_fp_add_23_8_0_cmp_3_b_core
      = bbox_req_stream_crt_sva_4_265_105[32:1];
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_4_inst_ccs_lp_piped_fp_add_23_8_0_cmp_4_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_4_inst_ccs_lp_piped_fp_add_23_8_0_cmp_4_b_core
      = bbox_req_stream_crt_sva_4_265_105[96:65];
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_5_inst_ccs_lp_piped_fp_add_23_8_0_cmp_5_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_5_inst_ccs_lp_piped_fp_add_23_8_0_cmp_5_b_core
      = bbox_req_stream_crt_sva_4_265_105[64:33];
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_6_inst_ccs_lp_piped_fp_add_23_8_0_cmp_6_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_6_inst_ccs_lp_piped_fp_add_23_8_0_cmp_6_b_core
      = bbox_req_stream_crt_sva_4_265_105[32:1];
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_7_inst_ccs_lp_piped_fp_add_23_8_0_cmp_7_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_7_inst_ccs_lp_piped_fp_add_23_8_0_cmp_7_b_core
      = bbox_req_stream_crt_sva_4_265_105[96:65];
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_8_inst_ccs_lp_piped_fp_add_23_8_0_cmp_8_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_8_inst_ccs_lp_piped_fp_add_23_8_0_cmp_8_b_core
      = bbox_req_stream_crt_sva_4_265_105[64:33];
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_9_inst_ccs_lp_piped_fp_add_23_8_0_cmp_9_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_9_inst_ccs_lp_piped_fp_add_23_8_0_cmp_9_b_core
      = bbox_req_stream_crt_sva_4_265_105[32:1];
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_10_inst_ccs_lp_piped_fp_add_23_8_0_cmp_10_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_10_inst_ccs_lp_piped_fp_add_23_8_0_cmp_10_b_core
      = bbox_req_stream_crt_sva_4_265_105[96:65];
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_11_inst_ccs_lp_piped_fp_add_23_8_0_cmp_11_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_11_inst_ccs_lp_piped_fp_add_23_8_0_cmp_11_b_core
      = bbox_req_stream_crt_sva_4_265_105[64:33];
  wire[7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_and_1_nl;
  wire[7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_if_acc_2_nl;
  wire[8:0] nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_if_acc_2_nl;
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_a_core;
  assign nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_if_acc_2_nl
      = conv_s2u_4_8({(leading_sign_8_0_1_0_out_3[3]) , (~ (leading_sign_8_0_1_0_out_3[2:0]))})
      + 8'b01111111;
  assign ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_if_acc_2_nl
      = nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_if_acc_2_nl[7:0];
  assign ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_and_1_nl
      = ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_if_acc_2_nl
      & (signext_8_1(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_x_u_sva_1[7]))
      & (signext_8_1(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_x_u_sva_1[7]));
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_a_core
      = {1'b0 , ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_and_1_nl
      , (ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_x_u_sva_1[6:0])
      , 16'b0000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_b_core
      = {1'b0 , (bbox_req_stream_rsci_idat_mxwt[273:266]) , 23'b00000000000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_1_a_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_1_a_core
      = bbox_req_stream_crt_sva_2_265_0[105:74];
  wire[7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_11_and_1_nl;
  wire[7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_11_if_acc_2_nl;
  wire[8:0] nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_11_if_acc_2_nl;
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_2_a_core;
  assign nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_11_if_acc_2_nl
      = conv_s2u_4_8({(leading_sign_8_0_1_0_11_out_3[3]) , (~ (leading_sign_8_0_1_0_11_out_3[2:0]))})
      + 8'b01111111;
  assign ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_11_if_acc_2_nl
      = nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_11_if_acc_2_nl[7:0];
  assign ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_11_and_1_nl
      = ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_11_if_acc_2_nl
      & (signext_8_1(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_11_x_u_sva_1[7]))
      & (signext_8_1(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_11_x_u_sva_1[7]));
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_2_a_core
      = {1'b0 , ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_11_and_1_nl
      , (ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_11_x_u_sva_1[6:0])
      , 16'b0000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_2_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_2_b_core
      = {1'b0 , (bbox_req_stream_rsci_idat_mxwt[289:282]) , 23'b00000000000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_3_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_3_a_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_3_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_3_a_core
      = bbox_req_stream_crt_sva_2_265_0[73:42];
  wire[7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_10_and_1_nl;
  wire[7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_10_if_acc_2_nl;
  wire[8:0] nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_10_if_acc_2_nl;
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_4_a_core;
  assign nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_10_if_acc_2_nl
      = conv_s2u_4_8({(leading_sign_8_0_1_0_10_out_3[3]) , (~ (leading_sign_8_0_1_0_10_out_3[2:0]))})
      + 8'b01111111;
  assign ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_10_if_acc_2_nl
      = nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_10_if_acc_2_nl[7:0];
  assign ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_10_and_1_nl
      = ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_10_if_acc_2_nl
      & (signext_8_1(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_10_x_u_sva_1[7]))
      & (signext_8_1(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_10_x_u_sva_1[7]));
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_4_a_core
      = {1'b0 , ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_10_and_1_nl
      , (ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_10_x_u_sva_1[6:0])
      , 16'b0000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_4_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_4_b_core
      = {1'b0 , (bbox_req_stream_rsci_idat_mxwt[281:274]) , 23'b00000000000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_5_a_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_5_a_core
      = bbox_req_stream_crt_sva_2_265_0[41:10];
  wire[7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_9_and_1_nl;
  wire[7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_9_if_acc_2_nl;
  wire[8:0] nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_9_if_acc_2_nl;
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_6_a_core;
  assign nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_9_if_acc_2_nl
      = conv_s2u_4_8({(leading_sign_8_0_1_0_9_out_3[3]) , (~ (leading_sign_8_0_1_0_9_out_3[2:0]))})
      + 8'b01111111;
  assign ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_9_if_acc_2_nl
      = nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_9_if_acc_2_nl[7:0];
  assign ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_9_and_1_nl
      = ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_9_if_acc_2_nl
      & (signext_8_1(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_9_x_u_sva_1[7]))
      & (signext_8_1(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_9_x_u_sva_1[7]));
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_6_a_core
      = {1'b0 , ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_9_and_1_nl
      , (ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_9_x_u_sva_1[6:0])
      , 16'b0000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_6_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_6_b_core
      = {1'b0 , (bbox_req_stream_rsci_idat_mxwt[273:266]) , 23'b00000000000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_7_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_7_a_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_7_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_7_a_core
      = bbox_req_stream_crt_sva_2_265_0[105:74];
  wire[7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_8_and_1_nl;
  wire[7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_8_if_acc_2_nl;
  wire[8:0] nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_8_if_acc_2_nl;
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_8_a_core;
  assign nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_8_if_acc_2_nl
      = conv_s2u_4_8({(leading_sign_8_0_1_0_8_out_3[3]) , (~ (leading_sign_8_0_1_0_8_out_3[2:0]))})
      + 8'b01111111;
  assign ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_8_if_acc_2_nl
      = nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_8_if_acc_2_nl[7:0];
  assign ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_8_and_1_nl
      = ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_8_if_acc_2_nl
      & (signext_8_1(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_8_x_u_sva_1[7]))
      & (signext_8_1(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_8_x_u_sva_1[7]));
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_8_a_core
      = {1'b0 , ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_8_and_1_nl
      , (ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_8_x_u_sva_1[6:0])
      , 16'b0000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_8_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_8_b_core
      = {1'b0 , (bbox_req_stream_rsci_idat_mxwt[289:282]) , 23'b00000000000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_9_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_9_a_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_9_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_9_a_core
      = bbox_req_stream_crt_sva_2_265_0[73:42];
  wire[7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_7_and_1_nl;
  wire[7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_7_if_acc_2_nl;
  wire[8:0] nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_7_if_acc_2_nl;
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_10_a_core;
  assign nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_7_if_acc_2_nl
      = conv_s2u_4_8({(leading_sign_8_0_1_0_7_out_3[3]) , (~ (leading_sign_8_0_1_0_7_out_3[2:0]))})
      + 8'b01111111;
  assign ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_7_if_acc_2_nl
      = nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_7_if_acc_2_nl[7:0];
  assign ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_7_and_1_nl
      = ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_7_if_acc_2_nl
      & (signext_8_1(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_7_x_u_sva_1[7]))
      & (signext_8_1(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_7_x_u_sva_1[7]));
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_10_a_core
      = {1'b0 , ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_7_and_1_nl
      , (ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_7_x_u_sva_1[6:0])
      , 16'b0000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_10_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_10_b_core
      = {1'b0 , (bbox_req_stream_rsci_idat_mxwt[281:274]) , 23'b00000000000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_11_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_11_a_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_11_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_11_a_core
      = bbox_req_stream_crt_sva_2_265_0[41:10];
  wire[7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_6_and_1_nl;
  wire[7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_6_if_acc_2_nl;
  wire[8:0] nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_6_if_acc_2_nl;
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_12_a_core;
  assign nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_6_if_acc_2_nl
      = conv_s2u_4_8({(leading_sign_8_0_1_0_6_out_3[3]) , (~ (leading_sign_8_0_1_0_6_out_3[2:0]))})
      + 8'b01111111;
  assign ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_6_if_acc_2_nl
      = nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_6_if_acc_2_nl[7:0];
  assign ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_6_and_1_nl
      = ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_6_if_acc_2_nl
      & (signext_8_1(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_6_x_u_sva_1[7]))
      & (signext_8_1(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_6_x_u_sva_1[7]));
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_12_a_core
      = {1'b0 , ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_6_and_1_nl
      , (ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_6_x_u_sva_1[6:0])
      , 16'b0000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_12_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_12_b_core
      = {1'b0 , (bbox_req_stream_rsci_idat_mxwt[273:266]) , 23'b00000000000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_13_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_13_a_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_13_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_13_a_core
      = bbox_req_stream_crt_sva_2_265_0[105:74];
  wire[7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_5_and_1_nl;
  wire[7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_5_if_acc_2_nl;
  wire[8:0] nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_5_if_acc_2_nl;
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_14_a_core;
  assign nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_5_if_acc_2_nl
      = conv_s2u_4_8({(leading_sign_8_0_1_0_5_out_3[3]) , (~ (leading_sign_8_0_1_0_5_out_3[2:0]))})
      + 8'b01111111;
  assign ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_5_if_acc_2_nl
      = nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_5_if_acc_2_nl[7:0];
  assign ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_5_and_1_nl
      = ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_5_if_acc_2_nl
      & (signext_8_1(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_5_x_u_sva_1[7]))
      & (signext_8_1(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_5_x_u_sva_1[7]));
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_14_a_core
      = {1'b0 , ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_5_and_1_nl
      , (ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_5_x_u_sva_1[6:0])
      , 16'b0000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_14_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_14_b_core
      = {1'b0 , (bbox_req_stream_rsci_idat_mxwt[289:282]) , 23'b00000000000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_15_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_15_a_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_15_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_15_a_core
      = bbox_req_stream_crt_sva_2_265_0[73:42];
  wire[7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_4_and_1_nl;
  wire[7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_4_if_acc_2_nl;
  wire[8:0] nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_4_if_acc_2_nl;
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_16_a_core;
  assign nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_4_if_acc_2_nl
      = conv_s2u_4_8({(leading_sign_8_0_1_0_4_out_3[3]) , (~ (leading_sign_8_0_1_0_4_out_3[2:0]))})
      + 8'b01111111;
  assign ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_4_if_acc_2_nl
      = nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_4_if_acc_2_nl[7:0];
  assign ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_4_and_1_nl
      = ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_4_if_acc_2_nl
      & (signext_8_1(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_4_x_u_sva_1[7]))
      & (signext_8_1(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_4_x_u_sva_1[7]));
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_16_a_core
      = {1'b0 , ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_4_and_1_nl
      , (ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_4_x_u_sva_1[6:0])
      , 16'b0000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_16_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_16_b_core
      = {1'b0 , (bbox_req_stream_rsci_idat_mxwt[281:274]) , 23'b00000000000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_17_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_17_a_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_17_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_17_a_core
      = bbox_req_stream_crt_sva_2_265_0[41:10];
  wire[7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_3_and_1_nl;
  wire[7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_3_if_acc_2_nl;
  wire[8:0] nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_3_if_acc_2_nl;
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_18_a_core;
  assign nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_3_if_acc_2_nl
      = conv_s2u_4_8({(leading_sign_8_0_1_0_3_out_3[3]) , (~ (leading_sign_8_0_1_0_3_out_3[2:0]))})
      + 8'b01111111;
  assign ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_3_if_acc_2_nl
      = nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_3_if_acc_2_nl[7:0];
  assign ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_3_and_1_nl
      = ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_3_if_acc_2_nl
      & (signext_8_1(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_3_x_u_sva_1[7]))
      & (signext_8_1(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_3_x_u_sva_1[7]));
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_18_a_core
      = {1'b0 , ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_3_and_1_nl
      , (ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_3_x_u_sva_1[6:0])
      , 16'b0000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_18_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_18_b_core
      = {1'b0 , (bbox_req_stream_rsci_idat_mxwt[273:266]) , 23'b00000000000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_19_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_19_a_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_19_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_19_a_core
      = bbox_req_stream_crt_sva_2_265_0[105:74];
  wire[7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_2_and_1_nl;
  wire[7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_2_if_acc_2_nl;
  wire[8:0] nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_2_if_acc_2_nl;
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_20_a_core;
  assign nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_2_if_acc_2_nl
      = conv_s2u_4_8({(leading_sign_8_0_1_0_2_out_3[3]) , (~ (leading_sign_8_0_1_0_2_out_3[2:0]))})
      + 8'b01111111;
  assign ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_2_if_acc_2_nl
      = nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_2_if_acc_2_nl[7:0];
  assign ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_2_and_1_nl
      = ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_2_if_acc_2_nl
      & (signext_8_1(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_2_x_u_sva_1[7]))
      & (signext_8_1(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_2_x_u_sva_1[7]));
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_20_a_core
      = {1'b0 , ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_2_and_1_nl
      , (ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_2_x_u_sva_1[6:0])
      , 16'b0000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_20_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_20_b_core
      = {1'b0 , (bbox_req_stream_rsci_idat_mxwt[289:282]) , 23'b00000000000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_21_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_21_a_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_21_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_21_a_core
      = bbox_req_stream_crt_sva_2_265_0[73:42];
  wire[7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_1_and_1_nl;
  wire[7:0] ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_1_if_acc_2_nl;
  wire[8:0] nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_1_if_acc_2_nl;
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_22_a_core;
  assign nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_1_if_acc_2_nl
      = conv_s2u_4_8({(leading_sign_8_0_1_0_1_out_3[3]) , (~ (leading_sign_8_0_1_0_1_out_3[2:0]))})
      + 8'b01111111;
  assign ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_1_if_acc_2_nl
      = nl_ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_1_if_acc_2_nl[7:0];
  assign ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_1_and_1_nl
      = ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_1_if_acc_2_nl
      & (signext_8_1(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_1_x_u_sva_1[7]))
      & (signext_8_1(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_1_x_u_sva_1[7]));
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_22_a_core
      = {1'b0 , ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_1_and_1_nl
      , (ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_1_x_u_sva_1[6:0])
      , 16'b0000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_22_b_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_22_b_core
      = {1'b0 , (bbox_req_stream_rsci_idat_mxwt[281:274]) , 23'b00000000000000000000000};
  wire [31:0] nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_23_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_23_a_core;
  assign nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_23_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_23_a_core
      = bbox_req_stream_crt_sva_2_265_0[41:10];
  wire  nl_bbox_core_staller_inst_core_flen_unreg;
  assign nl_bbox_core_staller_inst_core_flen_unreg = ~((~((~ and_17_tmp) & (fsm_output[1])))
      | and_211_cse | and_212_cse | and_213_cse | and_214_cse | and_215_cse | and_216_cse
      | and_217_cse | (main_stage_v_7 & (~(reg_bbox_resp_stream_rsci_iswt0_cse &
      (~ bbox_resp_stream_rsci_bawt))) & or_cse_1 & (fsm_output[1])) | (reg_bbox_resp_stream_rsci_iswt0_cse
      & or_cse_1 & (fsm_output[1])));
  ccs_dw_fp_cmp_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0)) ccs_fp_cmp_23_8_0_14_rg (
      .a(bbox_ns_fmax_return_d_2_lpi_1_dfm_1),
      .b(bbox_ns_fmax_return_d_5_lpi_1_dfm_1),
      .zctr(1'b0),
      .aeqb(ccs_fp_cmp_23_8_0_14_out_6),
      .altb(ccs_fp_cmp_23_8_0_14_out_7),
      .agtb(ccs_fp_cmp_23_8_0_14_out_8),
      .unordered(ccs_fp_cmp_23_8_0_14_out_9),
      .z0(ccs_fp_cmp_23_8_0_14_out_10),
      .z1(ccs_fp_cmp_23_8_0_14_out_11),
      .status0(status0_out),
      .status1(status1_out)
    );
  ccs_dw_fp_cmp_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0)) ccs_fp_cmp_23_8_0_13_rg (
      .a(bbox_ns_fmax_return_d_5_lpi_1_dfm_1),
      .b(return_ac_std_float_47_mux_itm_1),
      .zctr(1'b0),
      .aeqb(ccs_fp_cmp_23_8_0_13_out_6),
      .altb(ccs_fp_cmp_23_8_0_13_out_7),
      .agtb(ccs_fp_cmp_23_8_0_13_out_8),
      .unordered(ccs_fp_cmp_23_8_0_13_out_9),
      .z0(ccs_fp_cmp_23_8_0_13_out_10),
      .z1(ccs_fp_cmp_23_8_0_13_out_11),
      .status0(status0_out_1),
      .status1(status1_out_1)
    );
  ccs_dw_fp_cmp_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0)) ccs_fp_cmp_23_8_0_6_rg (
      .a(bbox_ns_fmax_return_d_2_lpi_1_dfm_1),
      .b(return_ac_std_float_23_mux_itm_1),
      .zctr(1'b0),
      .aeqb(ccs_fp_cmp_23_8_0_6_out_6),
      .altb(ccs_fp_cmp_23_8_0_6_out_7),
      .agtb(ccs_fp_cmp_23_8_0_6_out_8),
      .unordered(ccs_fp_cmp_23_8_0_6_out_9),
      .z0(ccs_fp_cmp_23_8_0_6_out_10),
      .z1(ccs_fp_cmp_23_8_0_6_out_11),
      .status0(status0_out_2),
      .status1(status1_out_2)
    );
  mgc_shift_l_v5 #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd8)) operator_8_false_11_lshift_rg (
      .a(bbox_ns_ldexpf_a_11_lpi_1_dfm_mx0),
      .s(leading_sign_8_0_1_0_11_out_3),
      .z(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_11_x_u_sva_1)
    );
  leading_sign_8_0_1_0  leading_sign_8_0_1_0_11_rg (
      .mantissa(bbox_ns_ldexpf_a_11_lpi_1_dfm_mx0),
      .rtn(leading_sign_8_0_1_0_11_out_3)
    );
  mgc_shift_l_v5 #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd8)) operator_8_false_10_lshift_rg (
      .a(bbox_ns_ldexpf_a_10_lpi_1_dfm_mx0),
      .s(leading_sign_8_0_1_0_10_out_3),
      .z(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_10_x_u_sva_1)
    );
  leading_sign_8_0_1_0  leading_sign_8_0_1_0_10_rg (
      .mantissa(bbox_ns_ldexpf_a_10_lpi_1_dfm_mx0),
      .rtn(leading_sign_8_0_1_0_10_out_3)
    );
  mgc_shift_l_v5 #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd8)) operator_8_false_9_lshift_rg (
      .a(bbox_ns_ldexpf_a_9_lpi_1_dfm_mx0),
      .s(leading_sign_8_0_1_0_9_out_3),
      .z(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_9_x_u_sva_1)
    );
  leading_sign_8_0_1_0  leading_sign_8_0_1_0_9_rg (
      .mantissa(bbox_ns_ldexpf_a_9_lpi_1_dfm_mx0),
      .rtn(leading_sign_8_0_1_0_9_out_3)
    );
  mgc_shift_l_v5 #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd8)) operator_8_false_8_lshift_rg (
      .a(bbox_ns_ldexpf_a_8_lpi_1_dfm_mx0),
      .s(leading_sign_8_0_1_0_8_out_3),
      .z(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_8_x_u_sva_1)
    );
  leading_sign_8_0_1_0  leading_sign_8_0_1_0_8_rg (
      .mantissa(bbox_ns_ldexpf_a_8_lpi_1_dfm_mx0),
      .rtn(leading_sign_8_0_1_0_8_out_3)
    );
  mgc_shift_l_v5 #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd8)) operator_8_false_7_lshift_rg (
      .a(bbox_ns_ldexpf_a_7_lpi_1_dfm_mx0),
      .s(leading_sign_8_0_1_0_7_out_3),
      .z(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_7_x_u_sva_1)
    );
  leading_sign_8_0_1_0  leading_sign_8_0_1_0_7_rg (
      .mantissa(bbox_ns_ldexpf_a_7_lpi_1_dfm_mx0),
      .rtn(leading_sign_8_0_1_0_7_out_3)
    );
  mgc_shift_l_v5 #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd8)) operator_8_false_6_lshift_rg (
      .a(bbox_ns_ldexpf_a_6_lpi_1_dfm_mx0),
      .s(leading_sign_8_0_1_0_6_out_3),
      .z(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_6_x_u_sva_1)
    );
  leading_sign_8_0_1_0  leading_sign_8_0_1_0_6_rg (
      .mantissa(bbox_ns_ldexpf_a_6_lpi_1_dfm_mx0),
      .rtn(leading_sign_8_0_1_0_6_out_3)
    );
  mgc_shift_l_v5 #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd8)) operator_8_false_5_lshift_rg (
      .a(bbox_ns_ldexpf_a_5_lpi_1_dfm_mx0),
      .s(leading_sign_8_0_1_0_5_out_3),
      .z(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_5_x_u_sva_1)
    );
  leading_sign_8_0_1_0  leading_sign_8_0_1_0_5_rg (
      .mantissa(bbox_ns_ldexpf_a_5_lpi_1_dfm_mx0),
      .rtn(leading_sign_8_0_1_0_5_out_3)
    );
  mgc_shift_l_v5 #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd8)) operator_8_false_4_lshift_rg (
      .a(bbox_ns_ldexpf_a_4_lpi_1_dfm_mx0),
      .s(leading_sign_8_0_1_0_4_out_3),
      .z(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_4_x_u_sva_1)
    );
  leading_sign_8_0_1_0  leading_sign_8_0_1_0_4_rg (
      .mantissa(bbox_ns_ldexpf_a_4_lpi_1_dfm_mx0),
      .rtn(leading_sign_8_0_1_0_4_out_3)
    );
  mgc_shift_l_v5 #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd8)) operator_8_false_3_lshift_rg (
      .a(bbox_ns_ldexpf_a_3_lpi_1_dfm_mx0),
      .s(leading_sign_8_0_1_0_3_out_3),
      .z(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_3_x_u_sva_1)
    );
  leading_sign_8_0_1_0  leading_sign_8_0_1_0_3_rg (
      .mantissa(bbox_ns_ldexpf_a_3_lpi_1_dfm_mx0),
      .rtn(leading_sign_8_0_1_0_3_out_3)
    );
  mgc_shift_l_v5 #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd8)) operator_8_false_2_lshift_rg (
      .a(bbox_ns_ldexpf_a_2_lpi_1_dfm_mx0),
      .s(leading_sign_8_0_1_0_2_out_3),
      .z(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_2_x_u_sva_1)
    );
  leading_sign_8_0_1_0  leading_sign_8_0_1_0_2_rg (
      .mantissa(bbox_ns_ldexpf_a_2_lpi_1_dfm_mx0),
      .rtn(leading_sign_8_0_1_0_2_out_3)
    );
  mgc_shift_l_v5 #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd8)) operator_8_false_1_lshift_rg (
      .a(bbox_ns_ldexpf_a_1_lpi_1_dfm_mx0),
      .s(leading_sign_8_0_1_0_1_out_3),
      .z(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_1_x_u_sva_1)
    );
  leading_sign_8_0_1_0  leading_sign_8_0_1_0_1_rg (
      .mantissa(bbox_ns_ldexpf_a_1_lpi_1_dfm_mx0),
      .rtn(leading_sign_8_0_1_0_1_out_3)
    );
  mgc_shift_l_v5 #(.width_a(32'sd8),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd8)) operator_8_false_lshift_rg (
      .a(bbox_ns_ldexpf_a_lpi_1_dfm_mx0),
      .s(leading_sign_8_0_1_0_out_3),
      .z(ac_std_float_cctor_assign_from_AC_RND_CONV_8_8_false_AC_TRN_AC_WRAP_x_u_sva_1)
    );
  leading_sign_8_0_1_0  leading_sign_8_0_1_0_rg (
      .mantissa(bbox_ns_ldexpf_a_lpi_1_dfm_mx0),
      .rtn(leading_sign_8_0_1_0_out_3)
    );
  ccs_dw_fp_cmp_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0)) ccs_fp_cmp_23_8_0_12_rg (
      .a(bbox_ns_fmin_return_d_3_lpi_1_dfm_mx0),
      .b(bbox_ns_fmin_return_d_4_lpi_1_dfm_mx0),
      .zctr(1'b0),
      .aeqb(ccs_fp_cmp_23_8_0_12_out_6),
      .altb(ccs_fp_cmp_23_8_0_12_out_7),
      .agtb(ccs_fp_cmp_23_8_0_12_out_8),
      .unordered(ccs_fp_cmp_23_8_0_12_out_9),
      .z0(ccs_fp_cmp_23_8_0_12_out_10),
      .z1(ccs_fp_cmp_23_8_0_12_out_11),
      .status0(status0_out_3),
      .status1(status1_out_3)
    );
  ccs_dw_fp_cmp_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0)) ccs_fp_cmp_23_8_0_11_rg (
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt),
      .b(nl_ccs_fp_cmp_23_8_0_11_rg_b[31:0]),
      .zctr(1'b0),
      .aeqb(ccs_fp_cmp_23_8_0_11_out_6),
      .altb(ccs_fp_cmp_23_8_0_11_out_7),
      .agtb(ccs_fp_cmp_23_8_0_11_out_8),
      .unordered(ccs_fp_cmp_23_8_0_11_out_9),
      .z0(ccs_fp_cmp_23_8_0_11_out_10),
      .z1(ccs_fp_cmp_23_8_0_11_out_11),
      .status0(status0_out_4),
      .status1(status1_out_4)
    );
  ccs_dw_fp_cmp_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0)) ccs_fp_cmp_23_8_0_10_rg (
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_3_z_mxwt),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt),
      .zctr(1'b0),
      .aeqb(ccs_fp_cmp_23_8_0_10_out_6),
      .altb(ccs_fp_cmp_23_8_0_10_out_7),
      .agtb(ccs_fp_cmp_23_8_0_10_out_8),
      .unordered(ccs_fp_cmp_23_8_0_10_out_9),
      .z0(ccs_fp_cmp_23_8_0_10_out_10),
      .z1(ccs_fp_cmp_23_8_0_10_out_11),
      .status0(status0_out_5),
      .status1(status1_out_5)
    );
  ccs_dw_fp_cmp_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0)) ccs_fp_cmp_23_8_0_9_rg (
      .a(bbox_ns_fmax_return_d_3_lpi_1_dfm_mx0),
      .b(bbox_ns_fmax_return_d_4_lpi_1_dfm_mx0),
      .zctr(1'b0),
      .aeqb(ccs_fp_cmp_23_8_0_9_out_6),
      .altb(ccs_fp_cmp_23_8_0_9_out_7),
      .agtb(ccs_fp_cmp_23_8_0_9_out_8),
      .unordered(ccs_fp_cmp_23_8_0_9_out_9),
      .z0(ccs_fp_cmp_23_8_0_9_out_10),
      .z1(ccs_fp_cmp_23_8_0_9_out_11),
      .status0(status0_out_6),
      .status1(status1_out_6)
    );
  ccs_dw_fp_cmp_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0)) ccs_fp_cmp_23_8_0_8_rg (
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_4_z_mxwt),
      .b(nl_ccs_fp_cmp_23_8_0_8_rg_b[31:0]),
      .zctr(1'b0),
      .aeqb(ccs_fp_cmp_23_8_0_8_out_6),
      .altb(ccs_fp_cmp_23_8_0_8_out_7),
      .agtb(ccs_fp_cmp_23_8_0_8_out_8),
      .unordered(ccs_fp_cmp_23_8_0_8_out_9),
      .z0(ccs_fp_cmp_23_8_0_8_out_10),
      .z1(ccs_fp_cmp_23_8_0_8_out_11),
      .status0(status0_out_7),
      .status1(status1_out_7)
    );
  ccs_dw_fp_cmp_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0)) ccs_fp_cmp_23_8_0_7_rg (
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_6_z_mxwt),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_5_z_mxwt),
      .zctr(1'b0),
      .aeqb(ccs_fp_cmp_23_8_0_7_out_6),
      .altb(ccs_fp_cmp_23_8_0_7_out_7),
      .agtb(ccs_fp_cmp_23_8_0_7_out_8),
      .unordered(ccs_fp_cmp_23_8_0_7_out_9),
      .z0(ccs_fp_cmp_23_8_0_7_out_10),
      .z1(ccs_fp_cmp_23_8_0_7_out_11),
      .status0(status0_out_8),
      .status1(status1_out_8)
    );
  ccs_dw_fp_cmp_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0)) ccs_fp_cmp_23_8_0_5_rg (
      .a(bbox_ns_fmin_return_d_lpi_1_dfm_mx0),
      .b(bbox_ns_fmin_return_d_1_lpi_1_dfm_mx0),
      .zctr(1'b0),
      .aeqb(ccs_fp_cmp_23_8_0_5_out_6),
      .altb(ccs_fp_cmp_23_8_0_5_out_7),
      .agtb(ccs_fp_cmp_23_8_0_5_out_8),
      .unordered(ccs_fp_cmp_23_8_0_5_out_9),
      .z0(ccs_fp_cmp_23_8_0_5_out_10),
      .z1(ccs_fp_cmp_23_8_0_5_out_11),
      .status0(status0_out_9),
      .status1(status1_out_9)
    );
  ccs_dw_fp_cmp_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0)) ccs_fp_cmp_23_8_0_4_rg (
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_7_z_mxwt),
      .b(nl_ccs_fp_cmp_23_8_0_4_rg_b[31:0]),
      .zctr(1'b0),
      .aeqb(ccs_fp_cmp_23_8_0_4_out_6),
      .altb(ccs_fp_cmp_23_8_0_4_out_7),
      .agtb(ccs_fp_cmp_23_8_0_4_out_8),
      .unordered(ccs_fp_cmp_23_8_0_4_out_9),
      .z0(ccs_fp_cmp_23_8_0_4_out_10),
      .z1(ccs_fp_cmp_23_8_0_4_out_11),
      .status0(status0_out_10),
      .status1(status1_out_10)
    );
  ccs_dw_fp_cmp_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0)) ccs_fp_cmp_23_8_0_3_rg (
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_9_z_mxwt),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_8_z_mxwt),
      .zctr(1'b0),
      .aeqb(ccs_fp_cmp_23_8_0_3_out_6),
      .altb(ccs_fp_cmp_23_8_0_3_out_7),
      .agtb(ccs_fp_cmp_23_8_0_3_out_8),
      .unordered(ccs_fp_cmp_23_8_0_3_out_9),
      .z0(ccs_fp_cmp_23_8_0_3_out_10),
      .z1(ccs_fp_cmp_23_8_0_3_out_11),
      .status0(status0_out_11),
      .status1(status1_out_11)
    );
  ccs_dw_fp_cmp_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0)) ccs_fp_cmp_23_8_0_2_rg (
      .a(bbox_ns_fmax_return_d_lpi_1_dfm_mx0),
      .b(bbox_ns_fmax_return_d_1_lpi_1_dfm_mx0),
      .zctr(1'b0),
      .aeqb(ccs_fp_cmp_23_8_0_2_out_6),
      .altb(ccs_fp_cmp_23_8_0_2_out_7),
      .agtb(ccs_fp_cmp_23_8_0_2_out_8),
      .unordered(ccs_fp_cmp_23_8_0_2_out_9),
      .z0(ccs_fp_cmp_23_8_0_2_out_10),
      .z1(ccs_fp_cmp_23_8_0_2_out_11),
      .status0(status0_out_12),
      .status1(status1_out_12)
    );
  ccs_dw_fp_cmp_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0)) ccs_fp_cmp_23_8_0_1_rg (
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_10_z_mxwt),
      .b(nl_ccs_fp_cmp_23_8_0_1_rg_b[31:0]),
      .zctr(1'b0),
      .aeqb(ccs_fp_cmp_23_8_0_1_out_6),
      .altb(ccs_fp_cmp_23_8_0_1_out_7),
      .agtb(ccs_fp_cmp_23_8_0_1_out_8),
      .unordered(ccs_fp_cmp_23_8_0_1_out_9),
      .z0(ccs_fp_cmp_23_8_0_1_out_10),
      .z1(ccs_fp_cmp_23_8_0_1_out_11),
      .status0(status0_out_13),
      .status1(status1_out_13)
    );
  ccs_dw_fp_cmp_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0)) ccs_fp_cmp_23_8_0_rg (
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt),
      .b(ccs_lp_piped_fp_add_23_8_0_cmp_11_z_mxwt),
      .zctr(1'b0),
      .aeqb(ccs_fp_cmp_23_8_0_out_6),
      .altb(ccs_fp_cmp_23_8_0_out_7),
      .agtb(ccs_fp_cmp_23_8_0_out_8),
      .unordered(ccs_fp_cmp_23_8_0_out_9),
      .z0(ccs_fp_cmp_23_8_0_out_10),
      .z1(ccs_fp_cmp_23_8_0_out_11),
      .status0(status0_out_14),
      .status1(status1_out_14)
    );
  bbox_core_bbox_req_stream_rsci bbox_core_bbox_req_stream_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .bbox_req_stream_rsc_dat(bbox_req_stream_rsc_dat),
      .bbox_req_stream_rsc_vld(bbox_req_stream_rsc_vld),
      .bbox_req_stream_rsc_rdy(bbox_req_stream_rsc_rdy),
      .core_wen(core_wen),
      .bbox_req_stream_rsci_oswt_unreg(and_211_cse),
      .bbox_req_stream_rsci_bawt(bbox_req_stream_rsci_bawt),
      .bbox_req_stream_rsci_iswt0(bbox_req_stream_rsci_iswt0),
      .bbox_req_stream_rsci_wen_comp(bbox_req_stream_rsci_wen_comp),
      .bbox_req_stream_rsci_idat_mxwt(bbox_req_stream_rsci_idat_mxwt)
    );
  bbox_core_bbox_resp_stream_rsci bbox_core_bbox_resp_stream_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .bbox_resp_stream_rsc_dat(bbox_resp_stream_rsc_dat),
      .bbox_resp_stream_rsc_vld(bbox_resp_stream_rsc_vld),
      .bbox_resp_stream_rsc_rdy(bbox_resp_stream_rsc_rdy),
      .core_wen(core_wen),
      .bbox_resp_stream_rsci_oswt_unreg(and_dcpl_6),
      .bbox_resp_stream_rsci_bawt(bbox_resp_stream_rsci_bawt),
      .bbox_resp_stream_rsci_iswt0(reg_bbox_resp_stream_rsci_iswt0_cse),
      .bbox_resp_stream_rsci_wen_comp(bbox_resp_stream_rsci_wen_comp),
      .bbox_resp_stream_rsci_idat(nl_bbox_core_bbox_resp_stream_rsci_inst_bbox_resp_stream_rsci_idat[204:0])
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_oswt_unreg(and_217_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_a_core(ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_b_core(nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_inst_ccs_lp_piped_fp_add_23_8_0_cmp_b_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_iswt1_pff(and_215_cse)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_1 bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_oswt_unreg(and_217_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_a_core(ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_b_core(nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_inst_ccs_lp_piped_fp_add_23_8_0_cmp_1_b_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1_pff(and_215_cse)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_2 bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_oswt_unreg(and_217_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_a_core(ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_b_core(nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_inst_ccs_lp_piped_fp_add_23_8_0_cmp_2_b_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1_pff(and_215_cse)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_3 bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_3_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_oswt_unreg(and_217_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_3_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_a_core(ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_b_core(nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_3_inst_ccs_lp_piped_fp_add_23_8_0_cmp_3_b_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_3_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1_pff(and_215_cse)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_4 bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_4_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_oswt_unreg(and_217_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_4_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_a_core(ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_b_core(nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_4_inst_ccs_lp_piped_fp_add_23_8_0_cmp_4_b_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_4_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1_pff(and_215_cse)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_5 bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_5_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_oswt_unreg(and_217_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_5_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_a_core(ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_b_core(nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_5_inst_ccs_lp_piped_fp_add_23_8_0_cmp_5_b_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_5_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1_pff(and_215_cse)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_6 bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_6_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_oswt_unreg(and_217_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_6_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_a_core(ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_b_core(nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_6_inst_ccs_lp_piped_fp_add_23_8_0_cmp_6_b_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_6_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1_pff(and_215_cse)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_7 bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_7_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_oswt_unreg(and_217_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_7_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_a_core(ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_b_core(nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_7_inst_ccs_lp_piped_fp_add_23_8_0_cmp_7_b_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_7_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1_pff(and_215_cse)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_8 bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_8_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_oswt_unreg(and_217_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_8_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_a_core(ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_b_core(nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_8_inst_ccs_lp_piped_fp_add_23_8_0_cmp_8_b_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_8_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1_pff(and_215_cse)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_9 bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_9_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_oswt_unreg(and_217_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_9_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_a_core(ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_b_core(nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_9_inst_ccs_lp_piped_fp_add_23_8_0_cmp_9_b_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_9_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1_pff(and_215_cse)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_10 bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_10_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_oswt_unreg(and_217_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_10_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_a_core(ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_b_core(nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_10_inst_ccs_lp_piped_fp_add_23_8_0_cmp_10_b_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_10_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1_pff(and_215_cse)
    );
  bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_11 bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_11_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_oswt_unreg(and_217_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_11_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_a_core(ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_b_core(nl_bbox_core_ccs_lp_piped_fp_add_23_8_0_cmp_11_inst_ccs_lp_piped_fp_add_23_8_0_cmp_11_b_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_11_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1_pff(and_215_cse)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_oswt_unreg(and_213_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_b_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1_pff(and_211_cse)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1 bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_oswt_unreg(and_215_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_1_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_b_core(ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1_pff(and_213_cse)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2 bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_oswt_unreg(and_213_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_2_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_b_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_2_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1_pff(and_211_cse)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_3 bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_3_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_oswt_unreg(and_215_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_3_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_3_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_3_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_b_core(ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1_pff(and_213_cse)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4 bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_oswt_unreg(and_213_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_4_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_b_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_4_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1_pff(and_211_cse)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5 bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_oswt_unreg(and_215_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_5_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_5_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_b_core(ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1_pff(and_213_cse)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6 bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_oswt_unreg(and_213_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_6_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_6_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_b_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_6_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1_pff(and_211_cse)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_7 bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_7_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_oswt_unreg(and_215_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_7_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_7_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_7_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_b_core(ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1_pff(and_213_cse)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8 bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_oswt_unreg(and_213_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_8_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_8_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_b_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_8_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1_pff(and_211_cse)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_9 bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_9_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_oswt_unreg(and_215_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_9_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_9_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_9_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_b_core(ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1_pff(and_213_cse)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10 bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_oswt_unreg(and_213_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_10_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_10_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_b_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_10_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1_pff(and_211_cse)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_11 bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_11_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_oswt_unreg(and_215_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_11_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_11_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_11_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_b_core(ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1_pff(and_213_cse)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12 bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_oswt_unreg(and_213_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_12_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_12_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_b_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_12_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1_pff(and_211_cse)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_13 bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_13_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_oswt_unreg(and_215_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_13_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_13_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_13_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_b_core(ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1_pff(and_213_cse)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14 bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_oswt_unreg(and_213_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_14_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_14_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_b_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_14_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1_pff(and_211_cse)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_15 bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_15_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_oswt_unreg(and_215_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_15_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_15_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_15_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_b_core(ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1_pff(and_213_cse)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16 bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_oswt_unreg(and_213_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_16_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_16_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_b_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_16_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1_pff(and_211_cse)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_17 bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_17_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_oswt_unreg(and_215_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_17_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_17_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_17_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_b_core(ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1_pff(and_213_cse)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18 bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_oswt_unreg(and_213_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_18_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_18_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_b_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_18_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1_pff(and_211_cse)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_19 bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_19_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_oswt_unreg(and_215_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_19_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_19_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_19_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_b_core(ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1_pff(and_213_cse)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20 bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_oswt_unreg(and_213_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_20_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_20_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_b_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_20_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1_pff(and_211_cse)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_21 bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_21_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_oswt_unreg(and_215_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_21_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_21_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_21_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_b_core(ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1_pff(and_213_cse)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22 bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_oswt_unreg(and_213_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_22_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_22_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_b_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_22_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1_pff(and_211_cse)
    );
  bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_23 bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_23_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_unreg(and_215_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_23_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_a_core(nl_bbox_core_ccs_lp_piped_fp_mult_23_8_0_cmp_23_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_23_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_b_core(ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1_pff(and_213_cse)
    );
  bbox_core_staller bbox_core_staller_inst (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .bbox_req_stream_rsci_wen_comp(bbox_req_stream_rsci_wen_comp),
      .bbox_resp_stream_rsci_wen_comp(bbox_resp_stream_rsci_wen_comp),
      .core_flen_unreg(nl_bbox_core_staller_inst_core_flen_unreg)
    );
  bbox_core_core_fsm bbox_core_core_fsm_inst (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign and_169_cse = core_wen & (~(reg_bbox_resp_stream_rsci_iswt0_cse & (~ bbox_resp_stream_rsci_bawt)))
      & main_stage_v_7;
  assign and_213_cse = and_13_tmp & (fsm_output[1]);
  assign and_215_cse = and_9_tmp & (fsm_output[1]);
  assign and_211_cse = and_17_tmp & (fsm_output[1]);
  assign and_217_cse = and_5_tmp & (fsm_output[1]);
  assign and_216_cse = and_7_tmp & (fsm_output[1]);
  assign and_214_cse = and_11_tmp & (fsm_output[1]);
  assign and_212_cse = and_15_tmp & (fsm_output[1]);
  assign bbox_req_stream_rid_and_1_cse = core_wen & and_5_tmp;
  assign and_187_cse = core_wen & (~((~ and_11_tmp) | (fsm_output[0])));
  assign and_192_cse = core_wen & (~((~ and_7_tmp) | (fsm_output[0])));
  assign and_197_cse = core_wen & (~((~ and_13_tmp) | (fsm_output[0])));
  assign and_199_cse = core_wen & (~((~ and_9_tmp) | (fsm_output[0])));
  assign and_17_tmp = bbox_req_stream_rsci_bawt & or_78_cse_1 & or_79_cse_1 & or_80_cse_1
      & or_81_cse_1 & or_82_cse_1 & or_83_cse_1 & or_84_cse_1 & or_85_cse_1 & or_86_cse_1
      & or_87_cse_1 & or_88_cse_1 & or_89_cse_1 & or_28_cse_1 & or_29_cse_1 & or_30_cse_1
      & or_31_cse_1 & or_32_cse_1 & or_33_cse_1 & or_34_cse_1 & or_35_cse_1 & or_36_cse_1
      & or_37_cse_1 & or_38_cse_1 & or_39_cse_1 & or_2_cse_1 & or_3_cse_1 & or_4_cse_1
      & or_5_cse_1 & or_6_cse_1 & or_7_cse_1 & or_8_cse_1 & or_9_cse_1 & or_10_cse_1
      & or_11_cse_1 & or_12_cse_1 & or_13_cse_1 & or_cse_1;
  assign and_15_tmp = main_stage_v_1 & or_78_cse_1 & or_79_cse_1 & or_80_cse_1 &
      or_81_cse_1 & or_82_cse_1 & or_83_cse_1 & or_84_cse_1 & or_85_cse_1 & or_86_cse_1
      & or_87_cse_1 & or_88_cse_1 & or_89_cse_1 & or_28_cse_1 & or_29_cse_1 & or_30_cse_1
      & or_31_cse_1 & or_32_cse_1 & or_33_cse_1 & or_34_cse_1 & or_35_cse_1 & or_36_cse_1
      & or_37_cse_1 & or_38_cse_1 & or_39_cse_1 & or_2_cse_1 & or_3_cse_1 & or_4_cse_1
      & or_5_cse_1 & or_6_cse_1 & or_7_cse_1 & or_8_cse_1 & or_9_cse_1 & or_10_cse_1
      & or_11_cse_1 & or_12_cse_1 & or_13_cse_1 & or_cse_1;
  assign and_13_tmp = main_stage_v_2 & or_78_cse_1 & or_79_cse_1 & or_80_cse_1 &
      or_81_cse_1 & or_82_cse_1 & or_83_cse_1 & or_84_cse_1 & or_85_cse_1 & or_86_cse_1
      & or_87_cse_1 & or_88_cse_1 & or_89_cse_1 & or_28_cse_1 & or_29_cse_1 & or_30_cse_1
      & or_31_cse_1 & or_32_cse_1 & or_33_cse_1 & or_34_cse_1 & or_35_cse_1 & or_36_cse_1
      & or_37_cse_1 & or_38_cse_1 & or_39_cse_1 & or_2_cse_1 & or_3_cse_1 & or_4_cse_1
      & or_5_cse_1 & or_6_cse_1 & or_7_cse_1 & or_8_cse_1 & or_9_cse_1 & or_10_cse_1
      & or_11_cse_1 & or_12_cse_1 & or_13_cse_1 & or_cse_1;
  assign and_11_tmp = main_stage_v_3 & or_28_cse_1 & or_29_cse_1 & or_30_cse_1 &
      or_31_cse_1 & or_32_cse_1 & or_33_cse_1 & or_34_cse_1 & or_35_cse_1 & or_36_cse_1
      & or_37_cse_1 & or_38_cse_1 & or_39_cse_1 & or_2_cse_1 & or_3_cse_1 & or_4_cse_1
      & or_5_cse_1 & or_6_cse_1 & or_7_cse_1 & or_8_cse_1 & or_9_cse_1 & or_10_cse_1
      & or_11_cse_1 & or_12_cse_1 & or_13_cse_1 & or_cse_1;
  assign and_9_tmp = main_stage_v_4 & or_28_cse_1 & or_29_cse_1 & or_30_cse_1 & or_31_cse_1
      & or_32_cse_1 & or_33_cse_1 & or_34_cse_1 & or_35_cse_1 & or_36_cse_1 & or_37_cse_1
      & or_38_cse_1 & or_39_cse_1 & or_2_cse_1 & or_3_cse_1 & or_4_cse_1 & or_5_cse_1
      & or_6_cse_1 & or_7_cse_1 & or_8_cse_1 & or_9_cse_1 & or_10_cse_1 & or_11_cse_1
      & or_12_cse_1 & or_13_cse_1 & or_cse_1;
  assign and_7_tmp = main_stage_v_5 & or_2_cse_1 & or_3_cse_1 & or_4_cse_1 & or_5_cse_1
      & or_6_cse_1 & or_7_cse_1 & or_8_cse_1 & or_9_cse_1 & or_10_cse_1 & or_11_cse_1
      & or_12_cse_1 & or_13_cse_1 & or_cse_1;
  assign and_5_tmp = main_stage_v_6 & or_2_cse_1 & or_3_cse_1 & or_4_cse_1 & or_5_cse_1
      & or_6_cse_1 & or_7_cse_1 & or_8_cse_1 & or_9_cse_1 & or_10_cse_1 & or_11_cse_1
      & or_12_cse_1 & or_13_cse_1 & or_cse_1;
  assign bbox_ns_ldexpf_a_11_lpi_1_dfm_mx0 = MUX_v_8_2_2((bbox_req_stream_rsci_idat_mxwt[385:378]),
      (bbox_req_stream_rsci_idat_mxwt[377:370]), bbox_req_stream_rsci_idat_mxwt[105]);
  assign bbox_ns_ldexpf_a_10_lpi_1_dfm_mx0 = MUX_v_8_2_2((bbox_req_stream_rsci_idat_mxwt[369:362]),
      (bbox_req_stream_rsci_idat_mxwt[361:354]), bbox_req_stream_rsci_idat_mxwt[73]);
  assign bbox_ns_ldexpf_a_9_lpi_1_dfm_mx0 = MUX_v_8_2_2((bbox_req_stream_rsci_idat_mxwt[353:346]),
      (bbox_req_stream_rsci_idat_mxwt[345:338]), bbox_req_stream_rsci_idat_mxwt[41]);
  assign bbox_ns_ldexpf_a_8_lpi_1_dfm_mx0 = MUX_v_8_2_2((bbox_req_stream_rsci_idat_mxwt[377:370]),
      (bbox_req_stream_rsci_idat_mxwt[385:378]), bbox_req_stream_rsci_idat_mxwt[105]);
  assign bbox_ns_ldexpf_a_7_lpi_1_dfm_mx0 = MUX_v_8_2_2((bbox_req_stream_rsci_idat_mxwt[361:354]),
      (bbox_req_stream_rsci_idat_mxwt[369:362]), bbox_req_stream_rsci_idat_mxwt[73]);
  assign bbox_ns_ldexpf_a_6_lpi_1_dfm_mx0 = MUX_v_8_2_2((bbox_req_stream_rsci_idat_mxwt[345:338]),
      (bbox_req_stream_rsci_idat_mxwt[353:346]), bbox_req_stream_rsci_idat_mxwt[41]);
  assign bbox_ns_ldexpf_a_5_lpi_1_dfm_mx0 = MUX_v_8_2_2((bbox_req_stream_rsci_idat_mxwt[337:330]),
      (bbox_req_stream_rsci_idat_mxwt[329:322]), bbox_req_stream_rsci_idat_mxwt[105]);
  assign bbox_ns_ldexpf_a_4_lpi_1_dfm_mx0 = MUX_v_8_2_2((bbox_req_stream_rsci_idat_mxwt[321:314]),
      (bbox_req_stream_rsci_idat_mxwt[313:306]), bbox_req_stream_rsci_idat_mxwt[73]);
  assign bbox_ns_ldexpf_a_3_lpi_1_dfm_mx0 = MUX_v_8_2_2((bbox_req_stream_rsci_idat_mxwt[305:298]),
      (bbox_req_stream_rsci_idat_mxwt[297:290]), bbox_req_stream_rsci_idat_mxwt[41]);
  assign bbox_ns_ldexpf_a_2_lpi_1_dfm_mx0 = MUX_v_8_2_2((bbox_req_stream_rsci_idat_mxwt[329:322]),
      (bbox_req_stream_rsci_idat_mxwt[337:330]), bbox_req_stream_rsci_idat_mxwt[105]);
  assign bbox_ns_ldexpf_a_1_lpi_1_dfm_mx0 = MUX_v_8_2_2((bbox_req_stream_rsci_idat_mxwt[313:306]),
      (bbox_req_stream_rsci_idat_mxwt[321:314]), bbox_req_stream_rsci_idat_mxwt[73]);
  assign bbox_ns_ldexpf_a_lpi_1_dfm_mx0 = MUX_v_8_2_2((bbox_req_stream_rsci_idat_mxwt[297:290]),
      (bbox_req_stream_rsci_idat_mxwt[305:298]), bbox_req_stream_rsci_idat_mxwt[41]);
  assign or_78_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_bawt | (~ main_stage_v_2);
  assign or_79_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_22_bawt | (~ main_stage_v_2);
  assign or_80_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_20_bawt | (~ main_stage_v_2);
  assign or_81_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_18_bawt | (~ main_stage_v_2);
  assign or_82_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_16_bawt | (~ main_stage_v_2);
  assign or_83_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_14_bawt | (~ main_stage_v_2);
  assign or_84_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_12_bawt | (~ main_stage_v_2);
  assign or_85_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_10_bawt | (~ main_stage_v_2);
  assign or_86_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_8_bawt | (~ main_stage_v_2);
  assign or_87_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_6_bawt | (~ main_stage_v_2);
  assign or_88_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt | (~ main_stage_v_2);
  assign or_89_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt | (~ main_stage_v_2);
  assign or_28_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_23_bawt | (~ main_stage_v_4);
  assign or_29_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_21_bawt | (~ main_stage_v_4);
  assign or_30_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_19_bawt | (~ main_stage_v_4);
  assign or_31_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_17_bawt | (~ main_stage_v_4);
  assign or_32_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_15_bawt | (~ main_stage_v_4);
  assign or_33_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_13_bawt | (~ main_stage_v_4);
  assign or_34_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_11_bawt | (~ main_stage_v_4);
  assign or_35_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_9_bawt | (~ main_stage_v_4);
  assign or_36_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_7_bawt | (~ main_stage_v_4);
  assign or_37_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_5_bawt | (~ main_stage_v_4);
  assign or_38_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_3_bawt | (~ main_stage_v_4);
  assign or_39_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt | (~ main_stage_v_4);
  assign or_2_cse_1 = ccs_lp_piped_fp_add_23_8_0_cmp_bawt | (~ main_stage_v_6);
  assign or_3_cse_1 = ccs_lp_piped_fp_add_23_8_0_cmp_11_bawt | (~ main_stage_v_6);
  assign or_4_cse_1 = ccs_lp_piped_fp_add_23_8_0_cmp_10_bawt | (~ main_stage_v_6);
  assign or_5_cse_1 = ccs_lp_piped_fp_add_23_8_0_cmp_9_bawt | (~ main_stage_v_6);
  assign or_6_cse_1 = ccs_lp_piped_fp_add_23_8_0_cmp_8_bawt | (~ main_stage_v_6);
  assign or_7_cse_1 = ccs_lp_piped_fp_add_23_8_0_cmp_7_bawt | (~ main_stage_v_6);
  assign or_8_cse_1 = ccs_lp_piped_fp_add_23_8_0_cmp_6_bawt | (~ main_stage_v_6);
  assign or_9_cse_1 = ccs_lp_piped_fp_add_23_8_0_cmp_5_bawt | (~ main_stage_v_6);
  assign or_10_cse_1 = ccs_lp_piped_fp_add_23_8_0_cmp_4_bawt | (~ main_stage_v_6);
  assign or_11_cse_1 = ccs_lp_piped_fp_add_23_8_0_cmp_3_bawt | (~ main_stage_v_6);
  assign or_12_cse_1 = ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt | (~ main_stage_v_6);
  assign or_13_cse_1 = ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt | (~ main_stage_v_6);
  assign or_cse_1 = bbox_resp_stream_rsci_bawt | (~ reg_bbox_resp_stream_rsci_iswt0_cse);
  assign FP_LEQ_32_8_11_nor_nl = ~(ccs_fp_cmp_23_8_0_11_out_7 | ccs_fp_cmp_23_8_0_11_out_6);
  assign bbox_ns_fmin_return_d_4_lpi_1_dfm_mx0 = MUX_v_32_2_2(ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt,
      (bbox_req_stream_crt_sva_6_265_202[63:32]), FP_LEQ_32_8_11_nor_nl);
  assign FP_LEQ_32_8_10_nor_nl = ~(ccs_fp_cmp_23_8_0_10_out_7 | ccs_fp_cmp_23_8_0_10_out_6);
  assign bbox_ns_fmin_return_d_3_lpi_1_dfm_mx0 = MUX_v_32_2_2(ccs_lp_piped_fp_add_23_8_0_cmp_3_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt, FP_LEQ_32_8_10_nor_nl);
  assign FP_LEQ_32_8_7_nor_nl = ~(ccs_fp_cmp_23_8_0_7_out_7 | ccs_fp_cmp_23_8_0_7_out_6);
  assign bbox_ns_fmax_return_d_3_lpi_1_dfm_mx0 = MUX_v_32_2_2(ccs_lp_piped_fp_add_23_8_0_cmp_5_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_6_z_mxwt, FP_LEQ_32_8_7_nor_nl);
  assign FP_LEQ_32_8_8_nor_nl = ~(ccs_fp_cmp_23_8_0_8_out_7 | ccs_fp_cmp_23_8_0_8_out_6);
  assign bbox_ns_fmax_return_d_4_lpi_1_dfm_mx0 = MUX_v_32_2_2((bbox_req_stream_crt_sva_6_265_202[31:0]),
      ccs_lp_piped_fp_add_23_8_0_cmp_4_z_mxwt, FP_LEQ_32_8_8_nor_nl);
  assign FP_LEQ_32_8_4_nor_nl = ~(ccs_fp_cmp_23_8_0_4_out_7 | ccs_fp_cmp_23_8_0_4_out_6);
  assign bbox_ns_fmin_return_d_1_lpi_1_dfm_mx0 = MUX_v_32_2_2(ccs_lp_piped_fp_add_23_8_0_cmp_7_z_mxwt,
      (bbox_req_stream_crt_sva_6_265_202[63:32]), FP_LEQ_32_8_4_nor_nl);
  assign FP_LEQ_32_8_3_nor_nl = ~(ccs_fp_cmp_23_8_0_3_out_7 | ccs_fp_cmp_23_8_0_3_out_6);
  assign bbox_ns_fmin_return_d_lpi_1_dfm_mx0 = MUX_v_32_2_2(ccs_lp_piped_fp_add_23_8_0_cmp_9_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_8_z_mxwt, FP_LEQ_32_8_3_nor_nl);
  assign FP_LEQ_32_8_nor_nl = ~(ccs_fp_cmp_23_8_0_out_7 | ccs_fp_cmp_23_8_0_out_6);
  assign bbox_ns_fmax_return_d_lpi_1_dfm_mx0 = MUX_v_32_2_2(ccs_lp_piped_fp_add_23_8_0_cmp_11_z_mxwt,
      ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt, FP_LEQ_32_8_nor_nl);
  assign FP_LEQ_32_8_1_nor_nl = ~(ccs_fp_cmp_23_8_0_1_out_7 | ccs_fp_cmp_23_8_0_1_out_6);
  assign bbox_ns_fmax_return_d_1_lpi_1_dfm_mx0 = MUX_v_32_2_2((bbox_req_stream_crt_sva_6_265_202[31:0]),
      ccs_lp_piped_fp_add_23_8_0_cmp_10_z_mxwt, FP_LEQ_32_8_1_nor_nl);
  assign and_dcpl_6 = reg_bbox_resp_stream_rsci_iswt0_cse & bbox_resp_stream_rsci_bawt;
  assign and_dcpl_7 = and_dcpl_6 & (~ main_stage_v_7);
  assign and_dcpl_12 = and_5_tmp & (~ bbox_req_stream_crt_sva_6_41);
  assign and_dcpl_14 = and_5_tmp & (~ bbox_req_stream_crt_sva_6_73);
  assign and_dcpl_16 = and_5_tmp & (~ bbox_req_stream_crt_sva_6_105);
  assign main_stage_v_7_mx0c1 = or_cse_1 & (~ and_5_tmp) & main_stage_v_7;
  assign main_stage_v_6_mx0c1 = and_5_tmp & (~ and_7_tmp) & (fsm_output[1]);
  assign main_stage_v_5_mx0c1 = and_7_tmp & (~ and_9_tmp) & (fsm_output[1]);
  assign main_stage_v_4_mx0c1 = and_9_tmp & (~ and_11_tmp) & (fsm_output[1]);
  assign main_stage_v_3_mx0c1 = and_11_tmp & (~ and_13_tmp) & (fsm_output[1]);
  assign main_stage_v_2_mx0c1 = and_13_tmp & (~ and_15_tmp) & (fsm_output[1]);
  assign main_stage_v_1_mx0c1 = and_15_tmp & (~ and_17_tmp) & (fsm_output[1]);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      bbox_req_stream_rsci_iswt0 <= 1'b0;
    end
    else if ( core_wen & (and_17_tmp | (fsm_output[0])) ) begin
      bbox_req_stream_rsci_iswt0 <= 1'b1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      bbox_resp_stream_rsci_idat_9_0 <= 10'b0000000000;
      bbox_resp_stream_rsci_idat_41_10 <= 32'b00000000000000000000000000000000;
      bbox_resp_stream_rsci_idat_73_42 <= 32'b00000000000000000000000000000000;
      bbox_resp_stream_rsci_idat_105_74 <= 32'b00000000000000000000000000000000;
      bbox_resp_stream_rsci_idat_137_106 <= 32'b00000000000000000000000000000000;
      bbox_resp_stream_rsci_idat_169_138 <= 32'b00000000000000000000000000000000;
      bbox_resp_stream_rsci_idat_201_170 <= 32'b00000000000000000000000000000000;
      bbox_resp_stream_rsci_idat_202 <= 1'b0;
      bbox_resp_stream_rsci_idat_203 <= 1'b0;
      bbox_resp_stream_rsci_idat_204 <= 1'b0;
    end
    else if ( and_169_cse ) begin
      bbox_resp_stream_rsci_idat_9_0 <= bbox_req_stream_rid_slc_bbox_req_stream_crt_9_0_itm_1;
      bbox_resp_stream_rsci_idat_41_10 <= const_x_min_ac_std_float_1_mux_itm_1;
      bbox_resp_stream_rsci_idat_73_42 <= const_z_min_ac_std_float_1_mux_itm_1;
      bbox_resp_stream_rsci_idat_105_74 <= const_z_min_ac_std_float_1_mux_1_itm_1;
      bbox_resp_stream_rsci_idat_137_106 <= const_x_min_ac_std_float_1_mux_1_itm_1;
      bbox_resp_stream_rsci_idat_169_138 <= const_z_min_ac_std_float_1_mux_2_itm_1;
      bbox_resp_stream_rsci_idat_201_170 <= const_z_min_ac_std_float_1_mux_3_itm_1;
      bbox_resp_stream_rsci_idat_202 <= ccs_fp_cmp_23_8_0_6_out_7 | ccs_fp_cmp_23_8_0_6_out_6;
      bbox_resp_stream_rsci_idat_203 <= ccs_fp_cmp_23_8_0_13_out_7 | ccs_fp_cmp_23_8_0_13_out_6;
      bbox_resp_stream_rsci_idat_204 <= ccs_fp_cmp_23_8_0_14_out_7 | ccs_fp_cmp_23_8_0_14_out_6;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1_cse <= 1'b0;
      reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_cse <= 1'b0;
      reg_ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1_cse <= 1'b0;
    end
    else if ( core_wen ) begin
      reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1_cse <= and_213_cse;
      reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_cse <= and_215_cse;
      reg_ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1_cse <= and_211_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_bbox_resp_stream_rsci_iswt0_cse <= 1'b0;
    end
    else if ( core_wen & ((or_cse_1 & main_stage_v_7) | and_dcpl_7) ) begin
      reg_bbox_resp_stream_rsci_iswt0_cse <= ~ and_dcpl_7;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_7 <= 1'b0;
    end
    else if ( core_wen & (and_217_cse | main_stage_v_7_mx0c1) ) begin
      main_stage_v_7 <= ~ main_stage_v_7_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      bbox_req_stream_rid_slc_bbox_req_stream_crt_9_0_itm_1 <= 10'b0000000000;
      const_x_min_ac_std_float_1_mux_itm_1 <= 32'b00000000000000000000000000000000;
      const_z_min_ac_std_float_1_mux_itm_1 <= 32'b00000000000000000000000000000000;
      const_z_min_ac_std_float_1_mux_3_itm_1 <= 32'b00000000000000000000000000000000;
      const_z_min_ac_std_float_1_mux_1_itm_1 <= 32'b00000000000000000000000000000000;
      const_z_min_ac_std_float_1_mux_2_itm_1 <= 32'b00000000000000000000000000000000;
      const_x_min_ac_std_float_1_mux_1_itm_1 <= 32'b00000000000000000000000000000000;
      bbox_ns_fmax_return_d_2_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      bbox_ns_fmax_return_d_5_lpi_1_dfm_1 <= 32'b00000000000000000000000000000000;
      return_ac_std_float_47_mux_itm_1 <= 32'b00000000000000000000000000000000;
      return_ac_std_float_23_mux_itm_1 <= 32'b00000000000000000000000000000000;
    end
    else if ( bbox_req_stream_rid_and_1_cse ) begin
      bbox_req_stream_rid_slc_bbox_req_stream_crt_9_0_itm_1 <= bbox_req_stream_crt_sva_6_9_0;
      const_x_min_ac_std_float_1_mux_itm_1 <= MUX_v_32_2_2(ccs_lp_piped_fp_add_23_8_0_cmp_9_z_mxwt,
          ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt, and_dcpl_12);
      const_z_min_ac_std_float_1_mux_itm_1 <= MUX_v_32_2_2(ccs_lp_piped_fp_add_23_8_0_cmp_8_z_mxwt,
          ccs_lp_piped_fp_add_23_8_0_cmp_11_z_mxwt, and_dcpl_14);
      const_z_min_ac_std_float_1_mux_3_itm_1 <= MUX_v_32_2_2(ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt,
          ccs_lp_piped_fp_add_23_8_0_cmp_4_z_mxwt, and_dcpl_16);
      const_z_min_ac_std_float_1_mux_1_itm_1 <= MUX_v_32_2_2(ccs_lp_piped_fp_add_23_8_0_cmp_7_z_mxwt,
          ccs_lp_piped_fp_add_23_8_0_cmp_10_z_mxwt, and_dcpl_16);
      const_z_min_ac_std_float_1_mux_2_itm_1 <= MUX_v_32_2_2(ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt,
          ccs_lp_piped_fp_add_23_8_0_cmp_5_z_mxwt, and_dcpl_14);
      const_x_min_ac_std_float_1_mux_1_itm_1 <= MUX_v_32_2_2(ccs_lp_piped_fp_add_23_8_0_cmp_3_z_mxwt,
          ccs_lp_piped_fp_add_23_8_0_cmp_6_z_mxwt, and_dcpl_12);
      bbox_ns_fmax_return_d_2_lpi_1_dfm_1 <= MUX_v_32_2_2(bbox_ns_fmax_return_d_1_lpi_1_dfm_mx0,
          bbox_ns_fmax_return_d_lpi_1_dfm_mx0, and_35_nl);
      bbox_ns_fmax_return_d_5_lpi_1_dfm_1 <= MUX_v_32_2_2(bbox_ns_fmax_return_d_4_lpi_1_dfm_mx0,
          bbox_ns_fmax_return_d_3_lpi_1_dfm_mx0, and_37_nl);
      return_ac_std_float_47_mux_itm_1 <= MUX_v_32_2_2(bbox_ns_fmin_return_d_3_lpi_1_dfm_mx0,
          bbox_ns_fmin_return_d_4_lpi_1_dfm_mx0, and_39_nl);
      return_ac_std_float_23_mux_itm_1 <= MUX_v_32_2_2(bbox_ns_fmin_return_d_lpi_1_dfm_mx0,
          bbox_ns_fmin_return_d_1_lpi_1_dfm_mx0, and_41_nl);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_6 <= 1'b0;
    end
    else if ( core_wen & (and_216_cse | main_stage_v_6_mx0c1) ) begin
      main_stage_v_6 <= ~ main_stage_v_6_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_5 <= 1'b0;
    end
    else if ( core_wen & (and_215_cse | main_stage_v_5_mx0c1) ) begin
      main_stage_v_5 <= ~ main_stage_v_5_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_4 <= 1'b0;
    end
    else if ( core_wen & (and_214_cse | main_stage_v_4_mx0c1) ) begin
      main_stage_v_4 <= ~ main_stage_v_4_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      bbox_req_stream_crt_sva_4_265_105 <= 161'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      bbox_req_stream_crt_sva_4_9_0 <= 10'b0000000000;
      bbox_req_stream_crt_sva_4_41 <= 1'b0;
      bbox_req_stream_crt_sva_4_73 <= 1'b0;
    end
    else if ( and_187_cse ) begin
      bbox_req_stream_crt_sva_4_265_105 <= bbox_req_stream_crt_sva_3_265_105;
      bbox_req_stream_crt_sva_4_9_0 <= bbox_req_stream_crt_sva_3_9_0;
      bbox_req_stream_crt_sva_4_41 <= bbox_req_stream_crt_sva_3_41;
      bbox_req_stream_crt_sva_4_73 <= bbox_req_stream_crt_sva_3_73;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_3 <= 1'b0;
    end
    else if ( core_wen & (and_213_cse | main_stage_v_3_mx0c1) ) begin
      main_stage_v_3 <= ~ main_stage_v_3_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_2 <= 1'b0;
    end
    else if ( core_wen & (and_212_cse | main_stage_v_2_mx0c1) ) begin
      main_stage_v_2 <= ~ main_stage_v_2_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      bbox_req_stream_crt_sva_2_265_0 <= 266'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ and_15_tmp) | (fsm_output[0]))) ) begin
      bbox_req_stream_crt_sva_2_265_0 <= bbox_req_stream_crt_sva_1_265_0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_1 <= 1'b0;
    end
    else if ( core_wen & (and_211_cse | main_stage_v_1_mx0c1) ) begin
      main_stage_v_1 <= ~ main_stage_v_1_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      bbox_req_stream_crt_sva_6_9_0 <= 10'b0000000000;
      bbox_req_stream_crt_sva_6_41 <= 1'b0;
      bbox_req_stream_crt_sva_6_73 <= 1'b0;
      bbox_req_stream_crt_sva_6_105 <= 1'b0;
      bbox_req_stream_crt_sva_6_265_202 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_192_cse ) begin
      bbox_req_stream_crt_sva_6_9_0 <= bbox_req_stream_crt_sva_5_9_0;
      bbox_req_stream_crt_sva_6_41 <= bbox_req_stream_crt_sva_5_41;
      bbox_req_stream_crt_sva_6_73 <= bbox_req_stream_crt_sva_5_73;
      bbox_req_stream_crt_sva_6_105 <= bbox_req_stream_crt_sva_5_105;
      bbox_req_stream_crt_sva_6_265_202 <= bbox_req_stream_crt_sva_5_265_202;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      bbox_req_stream_crt_sva_3_265_105 <= 161'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      bbox_req_stream_crt_sva_3_9_0 <= 10'b0000000000;
      bbox_req_stream_crt_sva_3_73 <= 1'b0;
      bbox_req_stream_crt_sva_3_41 <= 1'b0;
    end
    else if ( and_197_cse ) begin
      bbox_req_stream_crt_sva_3_265_105 <= bbox_req_stream_crt_sva_2_265_0[265:105];
      bbox_req_stream_crt_sva_3_9_0 <= bbox_req_stream_crt_sva_2_265_0[9:0];
      bbox_req_stream_crt_sva_3_73 <= bbox_req_stream_crt_sva_2_265_0[73];
      bbox_req_stream_crt_sva_3_41 <= bbox_req_stream_crt_sva_2_265_0[41];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      bbox_req_stream_crt_sva_1_265_0 <= 266'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( core_wen & (~((~ and_17_tmp) | (fsm_output[0]))) ) begin
      bbox_req_stream_crt_sva_1_265_0 <= bbox_req_stream_rsci_idat_mxwt[265:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      bbox_req_stream_crt_sva_5_265_202 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      bbox_req_stream_crt_sva_5_9_0 <= 10'b0000000000;
      bbox_req_stream_crt_sva_5_105 <= 1'b0;
      bbox_req_stream_crt_sva_5_41 <= 1'b0;
      bbox_req_stream_crt_sva_5_73 <= 1'b0;
    end
    else if ( and_199_cse ) begin
      bbox_req_stream_crt_sva_5_265_202 <= bbox_req_stream_crt_sva_4_265_105[160:97];
      bbox_req_stream_crt_sva_5_9_0 <= bbox_req_stream_crt_sva_4_9_0;
      bbox_req_stream_crt_sva_5_105 <= bbox_req_stream_crt_sva_4_265_105[0];
      bbox_req_stream_crt_sva_5_41 <= bbox_req_stream_crt_sva_4_41;
      bbox_req_stream_crt_sva_5_73 <= bbox_req_stream_crt_sva_4_73;
    end
  end
  assign and_35_nl = and_5_tmp & (~(ccs_fp_cmp_23_8_0_2_out_7 | ccs_fp_cmp_23_8_0_2_out_6));
  assign and_37_nl = and_5_tmp & (~(ccs_fp_cmp_23_8_0_9_out_7 | ccs_fp_cmp_23_8_0_9_out_6));
  assign and_39_nl = and_5_tmp & (~(ccs_fp_cmp_23_8_0_12_out_7 | ccs_fp_cmp_23_8_0_12_out_6));
  assign and_41_nl = and_5_tmp & (~(ccs_fp_cmp_23_8_0_5_out_7 | ccs_fp_cmp_23_8_0_5_out_6));

  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input  sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [7:0] signext_8_1;
    input  vector;
  begin
    signext_8_1= {{7{vector}}, vector};
  end
  endfunction


  function automatic [7:0] conv_s2u_4_8 ;
    input [3:0]  vector ;
  begin
    conv_s2u_4_8 = {{4{vector[3]}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist_core
// ------------------------------------------------------------------


module ist_core (
  clk, arst_n, ist_req_stream_rsc_dat, ist_req_stream_rsc_vld, ist_req_stream_rsc_rdy,
      ist_resp_stream_rsc_dat, ist_resp_stream_rsc_vld, ist_resp_stream_rsc_rdy
);
  input clk;
  input arst_n;
  input [553:0] ist_req_stream_rsc_dat;
  input ist_req_stream_rsc_vld;
  output ist_req_stream_rsc_rdy;
  output [106:0] ist_resp_stream_rsc_dat;
  output ist_resp_stream_rsc_vld;
  input ist_resp_stream_rsc_rdy;


  // Interconnect Declarations
  wire core_wen;
  wire core_wten;
  wire ist_req_stream_rsci_bawt;
  reg ist_req_stream_rsci_iswt0;
  wire ist_req_stream_rsci_wen_comp;
  wire [553:0] ist_req_stream_rsci_idat_mxwt;
  wire ist_resp_stream_rsci_bawt;
  wire ist_resp_stream_rsci_wen_comp;
  wire ccs_lp_piped_fp_recip_23_8_0_cmp_bawt;
  reg ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1;
  wire [31:0] ccs_lp_piped_fp_recip_23_8_0_cmp_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_3_bawt;
  reg ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_3_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_4_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_4_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_5_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_5_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_6_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_6_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_7_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_7_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_8_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_8_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_9_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_9_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_10_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_10_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_11_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_11_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_12_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_12_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_13_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_13_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_14_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_14_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_15_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_15_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_16_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_16_z_mxwt;
  wire ccs_lp_piped_fp_add_23_8_0_cmp_17_bawt;
  wire [31:0] ccs_lp_piped_fp_add_23_8_0_cmp_17_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_3_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt;
  reg ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_5_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_6_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_7_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_8_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_9_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_10_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_11_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_12_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_13_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_14_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_15_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_16_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_17_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_18_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_19_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_20_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_21_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_22_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_23_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_24_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_24_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_25_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_25_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_26_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_26_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_27_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_27_z_mxwt;
  wire ccs_lp_piped_fp_mult_23_8_0_cmp_28_bawt;
  wire [31:0] ccs_lp_piped_fp_mult_23_8_0_cmp_28_z_mxwt;
  reg [31:0] ist_resp_stream_rsci_idat_106_75;
  reg [31:0] ist_resp_stream_rsci_idat_74_43;
  reg [31:0] ist_resp_stream_rsci_idat_42_11;
  reg ist_resp_stream_rsci_idat_10;
  reg [9:0] ist_resp_stream_rsci_idat_9_0;
  reg ccs_lp_piped_fp_add_23_8_0_cmp_3_a_core_31;
  reg ccs_lp_piped_fp_add_23_8_0_cmp_3_b_core_31;
  wire [1:0] fsm_output;
  wire and_55_tmp;
  wire and_53_tmp;
  wire and_51_tmp;
  wire and_49_tmp;
  wire and_47_tmp;
  wire and_45_tmp;
  wire and_43_tmp;
  wire and_41_tmp;
  wire and_39_tmp;
  wire and_37_tmp;
  wire and_35_tmp;
  wire and_33_tmp;
  wire operator_1_false_1_xor_tmp;
  wire operator_1_false_xor_tmp;
  wire and_31_tmp;
  wire and_29_tmp;
  wire and_27_tmp;
  wire and_25_tmp;
  wire and_23_tmp;
  wire and_21_tmp;
  wire and_19_tmp;
  wire and_17_tmp;
  wire and_15_tmp;
  wire and_tmp;
  wire mux_tmp;
  wire and_tmp_1;
  wire nand_tmp_2;
  wire not_tmp_7;
  wire and_tmp_4;
  wire nor_tmp_15;
  wire mux_tmp_14;
  wire or_tmp_15;
  wire nand_tmp_3;
  wire mux_tmp_20;
  wire mux_tmp_21;
  wire mux_tmp_22;
  wire not_tmp_23;
  wire or_tmp_34;
  wire or_tmp_40;
  wire and_tmp_10;
  wire not_tmp_34;
  wire or_tmp_47;
  wire nand_tmp_11;
  wire mux_tmp_66;
  wire not_tmp_39;
  wire and_dcpl_4;
  wire and_dcpl_6;
  wire or_dcpl_5;
  wire and_dcpl_15;
  wire and_dcpl_20;
  wire and_dcpl_25;
  wire and_dcpl_37;
  wire and_dcpl_39;
  wire and_dcpl_40;
  wire and_dcpl_42;
  wire and_dcpl_47;
  wire or_dcpl_20;
  wire or_dcpl_25;
  wire and_dcpl_56;
  wire and_dcpl_61;
  wire or_dcpl_30;
  wire or_dcpl_34;
  wire and_dcpl_110;
  reg land_lpi_1_dfm_2;
  reg main_stage_v_21;
  wire or_523_cse_1;
  wire or_519_cse_1;
  wire or_1_cse_1;
  wire or_2_cse_1;
  wire or_3_cse_1;
  wire if_land_lpi_1_dfm_2;
  reg FP_GEQ_32_8_lor_lpi_1_dfm_2;
  reg main_stage_v_22;
  reg land_1_lpi_1_dfm_1_st_8;
  reg main_stage_v_23;
  reg main_stage_v_24;
  reg if_land_lpi_1_dfm_1_st_2;
  reg main_stage_v_25;
  reg main_stage_v_26;
  wire nand_5_cse_1;
  reg if_land_lpi_1_dfm_1_st_4;
  reg land_1_lpi_1_dfm_1_st_7;
  reg land_1_lpi_1_dfm_1_st_6;
  reg if_land_lpi_1_dfm_1_st_1;
  reg land_1_lpi_1_dfm_1_st_9;
  reg land_lpi_1_dfm_1;
  reg land_1_lpi_1_dfm_1_st_2;
  reg land_1_lpi_1_dfm_1_st_4;
  reg FP_LEQ_32_8_arelb_1_sva;
  reg fp_arelb_32_8_return_0_sva;
  reg [31:0] det_d_sva_2;
  wire and_632_cse;
  reg reg_ccs_lp_piped_fp_mult_23_8_0_cmp_28_iswt1_cse;
  reg reg_ccs_lp_piped_fp_mult_23_8_0_cmp_28_oswt_cse;
  reg reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_cse;
  reg reg_ccs_lp_piped_fp_mult_23_8_0_cmp_17_oswt_cse;
  reg reg_ccs_lp_piped_fp_mult_23_8_0_cmp_14_oswt_cse;
  reg reg_ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1_cse;
  reg reg_ccs_lp_piped_fp_mult_23_8_0_cmp_8_oswt_cse;
  reg reg_ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1_cse;
  reg reg_ccs_lp_piped_fp_add_23_8_0_cmp_8_oswt_cse;
  reg reg_ccs_lp_piped_fp_add_23_8_0_cmp_2_oswt_cse;
  wire det_d_and_cse;
  wire and_642_cse;
  wire if_aelse_and_2_cse;
  wire FP_LEQ_32_8_arelb_and_cse;
  wire aelse_and_cse;
  wire and_660_cse;
  wire det_d_and_4_cse;
  wire and_683_cse;
  wire det_d_and_3_cse;
  wire and_670_cse;
  wire det_d_and_7_cse;
  wire and_680_cse;
  wire and_673_cse;
  wire and_681_cse;
  wire aelse_1_and_4_cse;
  wire and_664_cse;
  wire aelse_1_and_11_cse;
  wire and_682_cse;
  wire aelse_1_and_5_cse;
  wire and_667_cse;
  wire aelse_1_and_12_cse;
  wire and_679_cse;
  wire aelse_1_and_6_cse;
  wire aelse_1_and_13_cse;
  wire aelse_and_2_cse;
  wire or_620_cse;
  wire and_751_cse;
  wire and_740_cse;
  wire nand_217_cse;
  wire or_561_cse;
  wire and_763_cse;
  wire and_761_cse;
  wire mux_151_cse;
  wire nand_223_cse;
  wire or_564_cse;
  wire or_607_cse;
  wire nand_228_cse;
  wire and_764_cse;
  reg reg_ist_resp_stream_rsci_iswt0_cse;
  wire and_776_cse;
  wire nand_206_cse;
  wire FP_LEQ_32_8_FP_LEQ_32_8_or_cse;
  wire lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_1_cse;
  wire lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_3_cse;
  wire lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_5_cse;
  wire lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_7_cse;
  wire lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_9_cse;
  wire lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_11_cse;
  wire lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_13_cse;
  wire lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_21_cse;
  wire lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_20_cse;
  wire lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_19_cse;
  wire lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_18_cse;
  wire lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_17_cse;
  wire lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_16_cse;
  wire lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_15_cse;
  wire lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_14_cse;
  wire lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_12_cse;
  wire lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_10_cse;
  wire lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_8_cse;
  wire lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_6_cse;
  wire lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_4_cse;
  wire lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_2_cse;
  wire nor_105_cse;
  wire and_744_cse;
  wire mux_131_cse;
  wire and_90_rmff;
  wire and_100_rmff;
  wire and_96_rmff;
  wire and_77_rmff;
  wire and_106_rmff;
  wire lp_piped_fp_add_AC_RND_CONV_0_32_8_15_mux1h_1_rmff;
  wire lp_piped_fp_add_AC_RND_CONV_0_32_8_15_mux1h_rmff;
  wire and_211_rmff;
  wire and_79_rmff;
  wire and_76_rmff;
  reg [31:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_23_sva_2;
  reg [31:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_20_sva_2;
  reg [31:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_17_sva_2;
  reg [31:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_14_sva_2;
  reg [31:0] ist_req_stream_crt_sva_20_265_234;
  reg [63:0] ist_req_stream_crt_sva_14_265_202;
  reg [31:0] c_z_d_sva_12;
  reg [31:0] n_z_d_sva_10;
  reg [31:0] c_y_d_sva_12;
  reg [31:0] n_y_d_sva_10;
  reg [31:0] c_x_d_sva_12;
  reg [31:0] n_x_d_sva_10;
  reg [191:0] ist_req_stream_crt_sva_6_553_362;
  reg [159:0] ist_req_stream_crt_sva_4_265_106;
  reg [30:0] det_d_sva_12_30_0;
  reg operator_1_false_return_1_sva_12;
  reg [30:0] vv_i_slc_vvv_d_30_0_itm_2;
  reg operator_1_false_return_sva_12;
  reg [30:0] uu_i_slc_uuu_d_30_0_itm_2;
  reg operator_1_false_return_2_sva_4;
  reg [30:0] if_tt_i_slc_if_ttt_d_30_0_itm_2;
  reg [31:0] det_d_sva_10;
  reg [31:0] det_d_sva_4;
  reg [159:0] ist_req_stream_crt_sva_2_265_106;
  wire [7:0] status0_out;
  wire [7:0] status1_out;
  wire [7:0] status0_out_1;
  wire [7:0] status1_out_1;
  wire [7:0] status0_out_2;
  wire [7:0] status1_out_2;
  reg main_stage_v_1;
  reg main_stage_v_2;
  reg main_stage_v_3;
  reg main_stage_v_4;
  reg main_stage_v_5;
  reg main_stage_v_6;
  reg main_stage_v_7;
  reg main_stage_v_8;
  reg main_stage_v_9;
  reg main_stage_v_10;
  reg main_stage_v_11;
  reg main_stage_v_12;
  reg main_stage_v_13;
  reg main_stage_v_14;
  reg main_stage_v_15;
  reg main_stage_v_16;
  reg main_stage_v_17;
  reg main_stage_v_18;
  reg main_stage_v_19;
  reg main_stage_v_20;
  reg FP_GEQ_32_8_lor_lpi_1_dfm_st;
  reg if_land_lpi_1_dfm_1_st;
  reg [31:0] n_x_d_sva_1;
  reg [31:0] n_x_d_sva_2;
  reg [31:0] n_x_d_sva_3;
  reg [31:0] n_x_d_sva_4;
  reg [31:0] n_x_d_sva_5;
  reg [31:0] n_x_d_sva_6;
  reg [31:0] n_x_d_sva_7;
  reg [31:0] n_x_d_sva_8;
  reg [31:0] n_x_d_sva_9;
  reg [31:0] n_y_d_sva_1;
  reg [31:0] n_y_d_sva_2;
  reg [31:0] n_y_d_sva_3;
  reg [31:0] n_y_d_sva_4;
  reg [31:0] n_y_d_sva_5;
  reg [31:0] n_y_d_sva_6;
  reg [31:0] n_y_d_sva_7;
  reg [31:0] n_y_d_sva_8;
  reg [31:0] n_y_d_sva_9;
  reg [31:0] n_z_d_sva_1;
  reg [31:0] n_z_d_sva_2;
  reg [31:0] n_z_d_sva_3;
  reg [31:0] n_z_d_sva_4;
  reg [31:0] n_z_d_sva_5;
  reg [31:0] n_z_d_sva_6;
  reg [31:0] n_z_d_sva_7;
  reg [31:0] n_z_d_sva_8;
  reg [31:0] n_z_d_sva_9;
  reg [31:0] c_x_d_sva_1;
  reg [31:0] c_x_d_sva_2;
  reg [31:0] c_x_d_sva_3;
  reg [31:0] c_x_d_sva_4;
  reg [31:0] c_x_d_sva_5;
  reg [31:0] c_x_d_sva_6;
  reg [31:0] c_x_d_sva_7;
  reg [31:0] c_x_d_sva_8;
  reg [31:0] c_x_d_sva_9;
  reg [31:0] c_x_d_sva_10;
  reg [31:0] c_x_d_sva_11;
  reg [31:0] c_y_d_sva_1;
  reg [31:0] c_y_d_sva_2;
  reg [31:0] c_y_d_sva_3;
  reg [31:0] c_y_d_sva_4;
  reg [31:0] c_y_d_sva_5;
  reg [31:0] c_y_d_sva_6;
  reg [31:0] c_y_d_sva_7;
  reg [31:0] c_y_d_sva_8;
  reg [31:0] c_y_d_sva_9;
  reg [31:0] c_y_d_sva_10;
  reg [31:0] c_y_d_sva_11;
  reg [31:0] c_z_d_sva_1;
  reg [31:0] c_z_d_sva_2;
  reg [31:0] c_z_d_sva_3;
  reg [31:0] c_z_d_sva_4;
  reg [31:0] c_z_d_sva_5;
  reg [31:0] c_z_d_sva_6;
  reg [31:0] c_z_d_sva_7;
  reg [31:0] c_z_d_sva_8;
  reg [31:0] c_z_d_sva_9;
  reg [31:0] c_z_d_sva_10;
  reg [31:0] c_z_d_sva_11;
  reg [31:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_14_sva_1;
  reg [31:0] det_d_sva_1;
  reg [31:0] det_d_sva_3;
  reg [31:0] det_d_sva_5;
  reg [31:0] det_d_sva_6;
  reg [31:0] det_d_sva_7;
  reg [31:0] det_d_sva_8;
  reg [31:0] det_d_sva_9;
  reg [31:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_17_sva_1;
  reg [31:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_20_sva_1;
  reg operator_1_false_return_sva_2;
  reg operator_1_false_return_sva_3;
  reg operator_1_false_return_sva_4;
  reg operator_1_false_return_sva_5;
  reg operator_1_false_return_sva_6;
  reg operator_1_false_return_sva_7;
  reg operator_1_false_return_sva_8;
  reg operator_1_false_return_sva_9;
  reg operator_1_false_return_sva_10;
  reg operator_1_false_return_sva_11;
  reg operator_1_false_return_1_sva_2;
  reg operator_1_false_return_1_sva_3;
  reg operator_1_false_return_1_sva_4;
  reg operator_1_false_return_1_sva_5;
  reg operator_1_false_return_1_sva_6;
  reg operator_1_false_return_1_sva_7;
  reg operator_1_false_return_1_sva_8;
  reg operator_1_false_return_1_sva_9;
  reg operator_1_false_return_1_sva_10;
  reg operator_1_false_return_1_sva_11;
  reg land_1_lpi_1_dfm_1_10;
  reg land_1_lpi_1_dfm_1_11;
  reg land_1_lpi_1_dfm_1_12;
  reg [31:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_23_sva_1;
  reg operator_1_false_return_2_sva_1;
  reg operator_1_false_return_2_sva_2;
  reg operator_1_false_return_2_sva_3;
  reg [31:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_24_sva_1;
  reg [31:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_24_sva_2;
  reg [31:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_24_sva_3;
  reg [31:0] lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_24_sva_4;
  reg if_land_lpi_1_dfm_1_3;
  reg [30:0] if_tt_i_slc_if_ttt_d_30_0_itm_1;
  reg [30:0] uu_i_slc_uuu_d_30_0_itm_1;
  reg [30:0] vv_i_slc_vvv_d_30_0_itm_1;
  reg if_if_if_if_and_itm_1;
  reg if_if_if_if_and_itm_2;
  reg if_if_if_if_and_itm_3;
  reg if_if_if_if_and_itm_4;
  reg [9:0] ist_req_stream_rid_slc_ist_req_stream_crt_9_0_itm_1;
  reg [9:0] ist_req_stream_rid_slc_ist_req_stream_crt_9_0_itm_2;
  reg [9:0] ist_req_stream_rid_slc_ist_req_stream_crt_9_0_itm_3;
  reg [9:0] ist_req_stream_rid_slc_ist_req_stream_crt_9_0_itm_4;
  reg [9:0] ist_req_stream_rid_slc_ist_req_stream_crt_9_0_itm_5;
  reg [9:0] ist_req_stream_rid_slc_ist_req_stream_crt_9_0_itm_6;
  reg land_1_lpi_1_dfm_1_st_1;
  reg land_1_lpi_1_dfm_1_st_3;
  reg land_1_lpi_1_dfm_1_st_5;
  reg [191:0] ist_req_stream_crt_sva_1_553_362;
  reg [159:0] ist_req_stream_crt_sva_1_265_106;
  reg [9:0] ist_req_stream_crt_sva_1_9_0;
  reg [191:0] ist_req_stream_crt_sva_2_553_362;
  reg [9:0] ist_req_stream_crt_sva_2_9_0;
  reg [191:0] ist_req_stream_crt_sva_3_553_362;
  reg [159:0] ist_req_stream_crt_sva_3_265_106;
  reg [9:0] ist_req_stream_crt_sva_3_9_0;
  reg [191:0] ist_req_stream_crt_sva_4_553_362;
  reg [9:0] ist_req_stream_crt_sva_4_9_0;
  reg [191:0] ist_req_stream_crt_sva_5_553_362;
  reg [63:0] ist_req_stream_crt_sva_5_265_202;
  reg [9:0] ist_req_stream_crt_sva_5_9_0;
  reg [63:0] ist_req_stream_crt_sva_6_265_202;
  reg [9:0] ist_req_stream_crt_sva_6_9_0;
  reg [63:0] ist_req_stream_crt_sva_7_265_202;
  reg [9:0] ist_req_stream_crt_sva_7_9_0;
  reg [63:0] ist_req_stream_crt_sva_8_265_202;
  reg [9:0] ist_req_stream_crt_sva_8_9_0;
  reg [63:0] ist_req_stream_crt_sva_9_265_202;
  reg [9:0] ist_req_stream_crt_sva_9_9_0;
  reg [63:0] ist_req_stream_crt_sva_10_265_202;
  reg [9:0] ist_req_stream_crt_sva_10_9_0;
  reg [63:0] ist_req_stream_crt_sva_11_265_202;
  reg [9:0] ist_req_stream_crt_sva_11_9_0;
  reg [63:0] ist_req_stream_crt_sva_12_265_202;
  reg [9:0] ist_req_stream_crt_sva_12_9_0;
  reg [63:0] ist_req_stream_crt_sva_13_265_202;
  reg [9:0] ist_req_stream_crt_sva_13_9_0;
  reg [9:0] ist_req_stream_crt_sva_14_9_0;
  reg [31:0] ist_req_stream_crt_sva_15_265_234;
  reg [9:0] ist_req_stream_crt_sva_15_9_0;
  reg [31:0] ist_req_stream_crt_sva_16_265_234;
  reg [9:0] ist_req_stream_crt_sva_16_9_0;
  reg [31:0] ist_req_stream_crt_sva_17_265_234;
  reg [9:0] ist_req_stream_crt_sva_17_9_0;
  reg [31:0] ist_req_stream_crt_sva_18_265_234;
  reg [9:0] ist_req_stream_crt_sva_18_9_0;
  reg [31:0] ist_req_stream_crt_sva_19_265_234;
  reg [9:0] ist_req_stream_crt_sva_19_9_0;
  reg [9:0] ist_req_stream_crt_sva_20_9_0;
  reg [30:0] det_d_sva_11_30_0;
  reg [30:0] uuu_d_sva_1_30_0;
  reg [30:0] uuu_d_sva_2_30_0;
  reg [30:0] uuu_d_sva_3_30_0;
  reg [30:0] uuu_d_sva_4_30_0;
  reg [30:0] uuu_d_sva_5_30_0;
  reg [30:0] uuu_d_sva_6_30_0;
  reg [30:0] uuu_d_sva_7_30_0;
  reg [30:0] uuu_d_sva_8_30_0;
  reg [30:0] uuu_d_sva_9_30_0;
  reg [30:0] uuu_d_sva_10_30_0;
  reg [30:0] vvv_d_sva_1_30_0;
  reg [30:0] vvv_d_sva_2_30_0;
  reg [30:0] vvv_d_sva_3_30_0;
  reg [30:0] vvv_d_sva_4_30_0;
  reg [30:0] vvv_d_sva_5_30_0;
  reg [30:0] vvv_d_sva_6_30_0;
  reg [30:0] vvv_d_sva_7_30_0;
  reg [30:0] vvv_d_sva_8_30_0;
  reg [30:0] vvv_d_sva_9_30_0;
  reg [30:0] vvv_d_sva_10_30_0;
  reg [30:0] if_ttt_d_sva_1_30_0;
  reg [30:0] if_ttt_d_sva_2_30_0;
  wire main_stage_v_21_mx0c1;
  wire main_stage_v_22_mx0c1;
  wire main_stage_v_23_mx0c1;
  wire main_stage_v_24_mx0c1;
  wire main_stage_v_25_mx0c1;
  wire main_stage_v_26_mx0c1;
  wire main_stage_v_20_mx0c1;
  wire main_stage_v_19_mx0c1;
  wire main_stage_v_18_mx0c1;
  wire main_stage_v_17_mx0c1;
  wire main_stage_v_16_mx0c1;
  wire main_stage_v_15_mx0c1;
  wire main_stage_v_14_mx0c1;
  wire main_stage_v_13_mx0c1;
  wire main_stage_v_12_mx0c1;
  wire main_stage_v_11_mx0c1;
  wire main_stage_v_10_mx0c1;
  wire main_stage_v_9_mx0c1;
  wire main_stage_v_8_mx0c1;
  wire main_stage_v_7_mx0c1;
  wire main_stage_v_6_mx0c1;
  wire main_stage_v_5_mx0c1;
  wire main_stage_v_4_mx0c1;
  wire main_stage_v_3_mx0c1;
  wire main_stage_v_2_mx0c1;
  wire main_stage_v_1_mx0c1;
  wire operator_1_false_return_2_sva_mx0w0;
  wire if_land_lpi_1_dfm_1_mx0w0;
  wire or_369_cse_1;
  wire or_370_cse_1;
  wire or_371_cse_1;
  wire or_372_cse_1;
  wire or_373_cse_1;
  wire or_374_cse_1;
  wire or_375_cse_1;
  wire or_376_cse_1;
  wire or_377_cse_1;
  wire or_289_cse_1;
  wire or_290_cse_1;
  wire or_291_cse_1;
  wire or_292_cse_1;
  wire or_293_cse_1;
  wire or_294_cse_1;
  wire or_295_cse_1;
  wire or_296_cse_1;
  wire or_297_cse_1;
  wire or_227_cse_1;
  wire or_228_cse_1;
  wire or_229_cse_1;
  wire or_230_cse_1;
  wire or_231_cse_1;
  wire or_232_cse_1;
  wire or_177_cse_1;
  wire or_178_cse_1;
  wire or_179_cse_1;
  wire or_180_cse_1;
  wire or_181_cse_1;
  wire or_182_cse_1;
  wire or_183_cse_1;
  wire or_141_cse_1;
  wire or_142_cse_1;
  wire or_143_cse_1;
  wire or_111_cse_1;
  wire or_112_cse_1;
  wire or_61_cse_1;
  wire or_62_cse_1;
  wire or_63_cse_1;
  wire or_64_cse_1;
  wire ccs_fp_cmp_23_8_0_2_out_6;
  wire ccs_fp_cmp_23_8_0_2_out_7;
  wire ccs_fp_cmp_23_8_0_2_out_8;
  wire ccs_fp_cmp_23_8_0_2_out_9;
  wire [31:0] ccs_fp_cmp_23_8_0_2_out_10;
  wire [31:0] ccs_fp_cmp_23_8_0_2_out_11;
  wire ccs_fp_cmp_23_8_0_1_out_6;
  wire ccs_fp_cmp_23_8_0_1_out_7;
  wire ccs_fp_cmp_23_8_0_1_out_8;
  wire ccs_fp_cmp_23_8_0_1_out_9;
  wire [31:0] ccs_fp_cmp_23_8_0_1_out_10;
  wire [31:0] ccs_fp_cmp_23_8_0_1_out_11;
  wire ccs_fp_cmp_23_8_0_out_6;
  wire ccs_fp_cmp_23_8_0_out_7;
  wire ccs_fp_cmp_23_8_0_out_8;
  wire ccs_fp_cmp_23_8_0_out_9;
  wire [31:0] ccs_fp_cmp_23_8_0_out_10;
  wire [31:0] ccs_fp_cmp_23_8_0_out_11;
  wire if_and_cse;
  wire and_799_cse;
  wire if_aelse_and_10_cse;
  wire and_801_cse;
  wire and_802_cse;
  wire if_ttt_d_and_2_cse;
  wire and_803_cse;
  wire aelse_1_and_26_cse;
  wire and_805_cse;
  wire and_806_cse;
  wire det_d_and_12_cse;
  wire aelse_1_and_28_cse;
  wire if_and_7_cse;
  wire det_d_and_15_cse;
  wire aelse_1_and_25_cse;
  wire if_and_10_cse;
  wire FP_GEQ_32_8_oelse_and_cse;
  wire and_815_cse;
  wire and_816_cse;
  wire and_743_cse;
  wire and_tmp_26;
  wire nand_245_cse;
  wire or_925_cse;
  wire or_924_cse;
  wire or_922_cse;
  wire or_920_cse;
  wire and_838_cse;

  wire mux_167_nl;
  wire and_850_nl;
  wire and_851_nl;
  wire mux_84_nl;
  wire and_58_nl;
  wire mux_83_nl;
  wire mux_82_nl;
  wire mux_79_nl;
  wire or_562_nl;
  wire mux_91_nl;
  wire mux_90_nl;
  wire mux_88_nl;
  wire or_570_nl;
  wire mux_87_nl;
  wire mux_86_nl;
  wire mux_85_nl;
  wire or_569_nl;
  wire mux_106_nl;
  wire and_765_nl;
  wire mux_105_nl;
  wire or_576_nl;
  wire mux_107_nl;
  wire and_767_nl;
  wire or_578_nl;
  wire mux_109_nl;
  wire and_771_nl;
  wire mux_108_nl;
  wire or_579_nl;
  wire mux_125_nl;
  wire mux_124_nl;
  wire mux_123_nl;
  wire mux_122_nl;
  wire mux_121_nl;
  wire mux_130_nl;
  wire and_780_nl;
  wire mux_129_nl;
  wire mux_128_nl;
  wire mux_127_nl;
  wire mux_126_nl;
  wire mux_138_nl;
  wire mux_136_nl;
  wire mux_166_nl;
  wire or_604_nl;
  wire and_787_nl;
  wire mux_143_nl;
  wire mux_142_nl;
  wire or_608_nl;
  wire mux_104_nl;
  wire mux_103_nl;
  wire mux_102_nl;
  wire mux_101_nl;
  wire mux_100_nl;
  wire mux_99_nl;
  wire or_575_nl;
  wire mux_98_nl;
  wire and_762_nl;
  wire mux_148_nl;
  wire and_791_nl;
  wire or_610_nl;
  wire nor_58_nl;
  wire or_581_nl;
  wire mux_78_nl;
  wire and_797_nl;
  wire mux_94_nl;
  wire mux_93_nl;
  wire mux_92_nl;
  wire nor_56_nl;
  wire mux_140_nl;
  wire mux_139_nl;
  wire mux_160_nl;
  wire nor_59_nl;
  wire mux_163_nl;
  wire or_656_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_ccs_fp_cmp_23_8_0_2_rg_a;
  assign nl_ccs_fp_cmp_23_8_0_2_rg_a = {operator_1_false_return_2_sva_2 , if_ttt_d_sva_2_30_0};
  wire [31:0] nl_ccs_fp_cmp_23_8_0_1_rg_a;
  assign nl_ccs_fp_cmp_23_8_0_1_rg_a = {operator_1_false_return_2_sva_mx0w0 , (ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt[30:0])};
  wire [31:0] nl_ccs_fp_cmp_23_8_0_rg_b;
  assign nl_ccs_fp_cmp_23_8_0_rg_b = {1'b0 , (det_d_sva_4[30:0])};
  wire [106:0] nl_ist_core_ist_resp_stream_rsci_inst_ist_resp_stream_rsci_idat;
  assign nl_ist_core_ist_resp_stream_rsci_inst_ist_resp_stream_rsci_idat = {ist_resp_stream_rsci_idat_106_75
      , ist_resp_stream_rsci_idat_74_43 , ist_resp_stream_rsci_idat_42_11 , ist_resp_stream_rsci_idat_10
      , ist_resp_stream_rsci_idat_9_0};
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_recip_23_8_0_cmp_inst_ccs_lp_piped_fp_recip_23_8_0_cmp_a_core;
  assign nl_ist_core_ccs_lp_piped_fp_recip_23_8_0_cmp_inst_ccs_lp_piped_fp_recip_23_8_0_cmp_a_core
      = {1'b0 , det_d_sva_12_30_0};
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_inst_ccs_lp_piped_fp_add_23_8_0_cmp_b_core;
  assign nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_inst_ccs_lp_piped_fp_add_23_8_0_cmp_b_core
      = {(~ (ccs_lp_piped_fp_mult_23_8_0_cmp_28_z_mxwt[31])) , (ccs_lp_piped_fp_mult_23_8_0_cmp_28_z_mxwt[30:0])};
  wire  nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_3_inst_ccs_lp_piped_fp_add_23_8_0_cmp_3_oswt_unreg;
  assign nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_3_inst_ccs_lp_piped_fp_add_23_8_0_cmp_3_oswt_unreg
      = land_lpi_1_dfm_2 & and_27_tmp;
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_3_inst_ccs_lp_piped_fp_add_23_8_0_cmp_3_a_core;
  assign nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_3_inst_ccs_lp_piped_fp_add_23_8_0_cmp_3_a_core
      = {lp_piped_fp_add_AC_RND_CONV_0_32_8_15_mux1h_1_rmff , (ccs_lp_piped_fp_add_23_8_0_cmp_6_z_mxwt[30:0])};
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_3_inst_ccs_lp_piped_fp_add_23_8_0_cmp_3_b_core;
  assign nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_3_inst_ccs_lp_piped_fp_add_23_8_0_cmp_3_b_core
      = {lp_piped_fp_add_AC_RND_CONV_0_32_8_15_mux1h_rmff , (ccs_lp_piped_fp_add_23_8_0_cmp_4_z_mxwt[30:0])};
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_10_inst_ccs_lp_piped_fp_add_23_8_0_cmp_10_b_core;
  assign nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_10_inst_ccs_lp_piped_fp_add_23_8_0_cmp_10_b_core
      = {(~ (ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_mxwt[31])) , (ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_mxwt[30:0])};
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_11_inst_ccs_lp_piped_fp_add_23_8_0_cmp_11_b_core;
  assign nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_11_inst_ccs_lp_piped_fp_add_23_8_0_cmp_11_b_core
      = {(~ (ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_mxwt[31])) , (ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_mxwt[30:0])};
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_12_inst_ccs_lp_piped_fp_add_23_8_0_cmp_12_b_core;
  assign nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_12_inst_ccs_lp_piped_fp_add_23_8_0_cmp_12_b_core
      = {(~ (ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_mxwt[31])) , (ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_mxwt[30:0])};
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_13_inst_ccs_lp_piped_fp_add_23_8_0_cmp_13_a_core;
  assign nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_13_inst_ccs_lp_piped_fp_add_23_8_0_cmp_13_a_core
      = ist_req_stream_rsci_idat_mxwt[361:330];
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_13_inst_ccs_lp_piped_fp_add_23_8_0_cmp_13_b_core;
  assign nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_13_inst_ccs_lp_piped_fp_add_23_8_0_cmp_13_b_core
      = {(~ (ist_req_stream_rsci_idat_mxwt[105])) , (ist_req_stream_rsci_idat_mxwt[104:74])};
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_14_inst_ccs_lp_piped_fp_add_23_8_0_cmp_14_a_core;
  assign nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_14_inst_ccs_lp_piped_fp_add_23_8_0_cmp_14_a_core
      = ist_req_stream_rsci_idat_mxwt[329:298];
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_14_inst_ccs_lp_piped_fp_add_23_8_0_cmp_14_b_core;
  assign nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_14_inst_ccs_lp_piped_fp_add_23_8_0_cmp_14_b_core
      = {(~ (ist_req_stream_rsci_idat_mxwt[73])) , (ist_req_stream_rsci_idat_mxwt[72:42])};
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_15_inst_ccs_lp_piped_fp_add_23_8_0_cmp_15_a_core;
  assign nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_15_inst_ccs_lp_piped_fp_add_23_8_0_cmp_15_a_core
      = ist_req_stream_rsci_idat_mxwt[297:266];
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_15_inst_ccs_lp_piped_fp_add_23_8_0_cmp_15_b_core;
  assign nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_15_inst_ccs_lp_piped_fp_add_23_8_0_cmp_15_b_core
      = {(~ (ist_req_stream_rsci_idat_mxwt[41])) , (ist_req_stream_rsci_idat_mxwt[40:10])};
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_16_inst_ccs_lp_piped_fp_add_23_8_0_cmp_16_b_core;
  assign nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_16_inst_ccs_lp_piped_fp_add_23_8_0_cmp_16_b_core
      = {(~ (ccs_lp_piped_fp_mult_23_8_0_cmp_24_z_mxwt[31])) , (ccs_lp_piped_fp_mult_23_8_0_cmp_24_z_mxwt[30:0])};
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_17_inst_ccs_lp_piped_fp_add_23_8_0_cmp_17_b_core;
  assign nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_17_inst_ccs_lp_piped_fp_add_23_8_0_cmp_17_b_core
      = {(~ (ccs_lp_piped_fp_mult_23_8_0_cmp_26_z_mxwt[31])) , (ccs_lp_piped_fp_mult_23_8_0_cmp_26_z_mxwt[30:0])};
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_a_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_a_core
      = ist_req_stream_rsci_idat_mxwt[425:394];
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_b_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_b_core
      = ist_req_stream_rsci_idat_mxwt[553:522];
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_1_b_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_1_b_core
      = {operator_1_false_return_1_sva_12 , vv_i_slc_vvv_d_30_0_itm_2};
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_2_b_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_2_b_core
      = {operator_1_false_return_sva_12 , uu_i_slc_uuu_d_30_0_itm_2};
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_3_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_3_b_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_3_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_3_b_core
      = {operator_1_false_return_2_sva_4 , if_tt_i_slc_if_ttt_d_30_0_itm_2};
  wire  nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_4_oswt_unreg;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_4_oswt_unreg
      = and_dcpl_15 & land_1_lpi_1_dfm_1_st_8 & ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt
      & FP_GEQ_32_8_lor_lpi_1_dfm_2 & main_stage_v_22;
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_4_a_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_4_a_core
      = {1'b0 , (det_d_sva_10[30:0])};
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_5_a_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_5_a_core
      = {1'b0 , (det_d_sva_4[30:0])};
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_5_b_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_5_b_core
      = ist_req_stream_crt_sva_14_265_202[31:0];
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_9_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_9_a_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_9_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_9_a_core
      = ist_req_stream_crt_sva_6_553_362[95:64];
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_10_a_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_10_a_core
      = ist_req_stream_crt_sva_6_553_362[63:32];
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_11_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_11_a_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_11_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_11_a_core
      = ist_req_stream_crt_sva_6_553_362[31:0];
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_12_a_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_12_a_core
      = ist_req_stream_crt_sva_6_553_362[191:160];
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_13_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_13_a_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_13_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_13_a_core
      = ist_req_stream_crt_sva_6_553_362[159:128];
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_14_a_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_14_a_core
      = ist_req_stream_crt_sva_6_553_362[127:96];
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_15_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_15_a_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_15_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_15_a_core
      = ist_req_stream_crt_sva_4_265_106[95:64];
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_16_a_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_16_a_core
      = ist_req_stream_crt_sva_4_265_106[63:32];
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_17_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_17_a_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_17_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_17_a_core
      = ist_req_stream_crt_sva_4_265_106[31:0];
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_18_a_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_18_a_core
      = ist_req_stream_crt_sva_2_265_106[63:32];
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_19_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_19_a_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_19_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_19_a_core
      = ist_req_stream_crt_sva_2_265_106[31:0];
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_20_a_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_20_a_core
      = ist_req_stream_crt_sva_2_265_106[31:0];
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_21_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_21_a_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_21_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_21_a_core
      = ist_req_stream_crt_sva_2_265_106[95:64];
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_22_a_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_22_a_core
      = ist_req_stream_crt_sva_2_265_106[95:64];
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_23_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_23_a_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_23_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_23_a_core
      = ist_req_stream_crt_sva_2_265_106[63:32];
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_24_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_24_a_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_24_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_24_a_core
      = ist_req_stream_rsci_idat_mxwt[425:394];
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_24_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_24_b_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_24_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_24_b_core
      = ist_req_stream_rsci_idat_mxwt[489:458];
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_25_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_25_a_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_25_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_25_a_core
      = ist_req_stream_rsci_idat_mxwt[393:362];
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_25_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_25_b_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_25_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_25_b_core
      = ist_req_stream_rsci_idat_mxwt[521:490];
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_26_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_26_a_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_26_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_26_a_core
      = ist_req_stream_rsci_idat_mxwt[393:362];
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_26_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_26_b_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_26_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_26_b_core
      = ist_req_stream_rsci_idat_mxwt[553:522];
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_27_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_27_a_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_27_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_27_a_core
      = ist_req_stream_rsci_idat_mxwt[457:426];
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_27_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_27_b_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_27_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_27_b_core
      = ist_req_stream_rsci_idat_mxwt[489:458];
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_28_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_28_a_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_28_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_28_a_core
      = ist_req_stream_rsci_idat_mxwt[457:426];
  wire [31:0] nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_28_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_28_b_core;
  assign nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_28_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_28_b_core
      = ist_req_stream_rsci_idat_mxwt[521:490];
  wire  nl_ist_core_staller_inst_core_flen_unreg;
  assign nl_ist_core_staller_inst_core_flen_unreg = ~((~((~ and_55_tmp) & (fsm_output[1])))
      | lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_1_cse
      | lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_2_cse
      | lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_3_cse
      | lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_4_cse
      | lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_5_cse
      | lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_6_cse
      | lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_7_cse
      | lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_8_cse
      | lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_9_cse
      | lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_10_cse
      | lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_11_cse
      | lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_12_cse
      | lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_13_cse
      | lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_14_cse
      | lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_15_cse
      | lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_16_cse
      | lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_17_cse
      | lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_18_cse
      | lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_19_cse
      | lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_20_cse
      | lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_21_cse
      | (main_stage_v_21 & (~(main_stage_v_22 & (or_dcpl_20 | (land_1_lpi_1_dfm_1_st_8
      & (~ ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt) & FP_GEQ_32_8_lor_lpi_1_dfm_2))))
      & or_523_cse_1 & or_519_cse_1 & or_1_cse_1 & or_2_cse_1 & or_3_cse_1 & or_925_cse
      & (fsm_output[1])) | (main_stage_v_22 & (~(main_stage_v_23 & or_dcpl_25)) &
      or_523_cse_1 & or_519_cse_1 & or_1_cse_1 & or_2_cse_1 & or_3_cse_1 & or_925_cse
      & (fsm_output[1])) | (main_stage_v_23 & (~(main_stage_v_24 & (or_dcpl_30 |
      ((~ ccs_lp_piped_fp_recip_23_8_0_cmp_bawt) & if_land_lpi_1_dfm_1_st_2 & land_1_lpi_1_dfm_1_10))))
      & or_519_cse_1 & or_1_cse_1 & or_2_cse_1 & or_3_cse_1 & or_925_cse & (fsm_output[1]))
      | (main_stage_v_24 & (~(main_stage_v_25 & or_dcpl_34)) & or_519_cse_1 & or_1_cse_1
      & or_2_cse_1 & or_3_cse_1 & or_925_cse & (fsm_output[1])) | (main_stage_v_25
      & (~(main_stage_v_26 & or_dcpl_5)) & or_1_cse_1 & or_2_cse_1 & or_3_cse_1 &
      or_925_cse & (fsm_output[1])) | (main_stage_v_26 & (~(reg_ist_resp_stream_rsci_iswt0_cse
      & (~ ist_resp_stream_rsci_bawt))) & or_1_cse_1 & or_2_cse_1 & or_3_cse_1 &
      or_925_cse & (fsm_output[1])) | (reg_ist_resp_stream_rsci_iswt0_cse & or_925_cse
      & (fsm_output[1])));
  ccs_dw_fp_cmp_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0)) ccs_fp_cmp_23_8_0_2_rg (
      .a(nl_ccs_fp_cmp_23_8_0_2_rg_a[31:0]),
      .b(ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_mxwt),
      .zctr(1'b0),
      .aeqb(ccs_fp_cmp_23_8_0_2_out_6),
      .altb(ccs_fp_cmp_23_8_0_2_out_7),
      .agtb(ccs_fp_cmp_23_8_0_2_out_8),
      .unordered(ccs_fp_cmp_23_8_0_2_out_9),
      .z0(ccs_fp_cmp_23_8_0_2_out_10),
      .z1(ccs_fp_cmp_23_8_0_2_out_11),
      .status0(status0_out),
      .status1(status1_out)
    );
  ccs_dw_fp_cmp_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0)) ccs_fp_cmp_23_8_0_1_rg (
      .a(nl_ccs_fp_cmp_23_8_0_1_rg_a[31:0]),
      .b(lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_24_sva_4),
      .zctr(1'b0),
      .aeqb(ccs_fp_cmp_23_8_0_1_out_6),
      .altb(ccs_fp_cmp_23_8_0_1_out_7),
      .agtb(ccs_fp_cmp_23_8_0_1_out_8),
      .unordered(ccs_fp_cmp_23_8_0_1_out_9),
      .z0(ccs_fp_cmp_23_8_0_1_out_10),
      .z1(ccs_fp_cmp_23_8_0_1_out_11),
      .status0(status0_out_1),
      .status1(status1_out_1)
    );
  ccs_dw_fp_cmp_v1 #(.sig_width(32'sd23),
  .exp_width(32'sd8),
  .ieee_compliance(32'sd0)) ccs_fp_cmp_23_8_0_rg (
      .a(ccs_lp_piped_fp_add_23_8_0_cmp_3_z_mxwt),
      .b(nl_ccs_fp_cmp_23_8_0_rg_b[31:0]),
      .zctr(1'b0),
      .aeqb(ccs_fp_cmp_23_8_0_out_6),
      .altb(ccs_fp_cmp_23_8_0_out_7),
      .agtb(ccs_fp_cmp_23_8_0_out_8),
      .unordered(ccs_fp_cmp_23_8_0_out_9),
      .z0(ccs_fp_cmp_23_8_0_out_10),
      .z1(ccs_fp_cmp_23_8_0_out_11),
      .status0(status0_out_2),
      .status1(status1_out_2)
    );
  ist_core_ist_req_stream_rsci ist_core_ist_req_stream_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .ist_req_stream_rsc_dat(ist_req_stream_rsc_dat),
      .ist_req_stream_rsc_vld(ist_req_stream_rsc_vld),
      .ist_req_stream_rsc_rdy(ist_req_stream_rsc_rdy),
      .core_wen(core_wen),
      .ist_req_stream_rsci_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_1_cse),
      .ist_req_stream_rsci_bawt(ist_req_stream_rsci_bawt),
      .ist_req_stream_rsci_iswt0(ist_req_stream_rsci_iswt0),
      .ist_req_stream_rsci_wen_comp(ist_req_stream_rsci_wen_comp),
      .ist_req_stream_rsci_idat_mxwt(ist_req_stream_rsci_idat_mxwt)
    );
  ist_core_ist_resp_stream_rsci ist_core_ist_resp_stream_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .ist_resp_stream_rsc_dat(ist_resp_stream_rsc_dat),
      .ist_resp_stream_rsc_vld(ist_resp_stream_rsc_vld),
      .ist_resp_stream_rsc_rdy(ist_resp_stream_rsc_rdy),
      .core_wen(core_wen),
      .ist_resp_stream_rsci_oswt_unreg(and_dcpl_39),
      .ist_resp_stream_rsci_bawt(ist_resp_stream_rsci_bawt),
      .ist_resp_stream_rsci_iswt0(reg_ist_resp_stream_rsci_iswt0_cse),
      .ist_resp_stream_rsci_wen_comp(ist_resp_stream_rsci_wen_comp),
      .ist_resp_stream_rsci_idat(nl_ist_core_ist_resp_stream_rsci_inst_ist_resp_stream_rsci_idat[106:0])
    );
  ist_core_ccs_lp_piped_fp_recip_23_8_0_cmp ist_core_ccs_lp_piped_fp_recip_23_8_0_cmp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_oswt_unreg(and_90_rmff),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_bawt(ccs_lp_piped_fp_recip_23_8_0_cmp_bawt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1(ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_a_core(nl_ist_core_ccs_lp_piped_fp_recip_23_8_0_cmp_inst_ccs_lp_piped_fp_recip_23_8_0_cmp_a_core[31:0]),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_z_mxwt(ccs_lp_piped_fp_recip_23_8_0_cmp_z_mxwt),
      .ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1_pff(and_106_rmff)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_5_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_28_oswt_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_a_core(ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_b_core(nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_inst_ccs_lp_piped_fp_add_23_8_0_cmp_b_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_3_cse)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_1 ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_oswt_unreg(and_764_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1(reg_ccs_lp_piped_fp_add_23_8_0_cmp_2_oswt_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_a_core(ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_b_core(lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_23_sva_2),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_1_iswt1_pff(and_100_rmff)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_2 ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_2_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_oswt_unreg(and_100_rmff),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_8_oswt_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_a_core(ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_b_core(ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_2_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_2_iswt1_pff(and_77_rmff)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_3 ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_3_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_oswt_unreg(nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_3_inst_ccs_lp_piped_fp_add_23_8_0_cmp_3_oswt_unreg),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_3_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1(ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_a_core(nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_3_inst_ccs_lp_piped_fp_add_23_8_0_cmp_3_a_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_b_core(nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_3_inst_ccs_lp_piped_fp_add_23_8_0_cmp_3_b_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_3_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1_pff(and_211_rmff)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_4 ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_4_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_13_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_4_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1(reg_ccs_lp_piped_fp_add_23_8_0_cmp_8_oswt_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_a_core(ccs_lp_piped_fp_add_23_8_0_cmp_5_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_b_core(lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_20_sva_2),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_4_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_4_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_11_cse)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_5 ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_5_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_11_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_5_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_14_oswt_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_a_core(ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_b_core(ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_5_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_5_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_9_cse)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_6 ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_6_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_13_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_6_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1(reg_ccs_lp_piped_fp_add_23_8_0_cmp_8_oswt_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_a_core(ccs_lp_piped_fp_add_23_8_0_cmp_7_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_b_core(lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_17_sva_2),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_6_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_6_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_11_cse)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_7 ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_7_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_11_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_7_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_14_oswt_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_a_core(ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_b_core(ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_7_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_7_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_9_cse)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_8 ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_8_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_11_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_8_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_14_oswt_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_a_core(ccs_lp_piped_fp_add_23_8_0_cmp_9_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_b_core(lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_14_sva_2),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_8_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_8_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_9_cse)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_9 ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_9_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_9_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_9_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_17_oswt_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_a_core(ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_b_core(ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_9_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_9_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_7_cse)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_10 ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_10_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_7_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_10_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_a_core(ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_b_core(nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_10_inst_ccs_lp_piped_fp_add_23_8_0_cmp_10_b_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_10_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_10_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_5_cse)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_11 ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_11_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_7_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_11_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_a_core(ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_b_core(nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_11_inst_ccs_lp_piped_fp_add_23_8_0_cmp_11_b_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_11_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_11_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_5_cse)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_12 ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_12_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_12_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_7_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_12_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_12_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_12_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_12_a_core(ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_12_b_core(nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_12_inst_ccs_lp_piped_fp_add_23_8_0_cmp_12_b_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_12_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_12_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_12_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_5_cse)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_13 ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_13_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_13_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_3_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_13_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_13_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_13_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_28_iswt1_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_13_a_core(nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_13_inst_ccs_lp_piped_fp_add_23_8_0_cmp_13_a_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_13_b_core(nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_13_inst_ccs_lp_piped_fp_add_23_8_0_cmp_13_b_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_13_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_13_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_13_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_1_cse)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_14 ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_14_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_14_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_3_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_14_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_14_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_14_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_28_iswt1_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_14_a_core(nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_14_inst_ccs_lp_piped_fp_add_23_8_0_cmp_14_a_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_14_b_core(nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_14_inst_ccs_lp_piped_fp_add_23_8_0_cmp_14_b_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_14_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_14_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_14_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_1_cse)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_15 ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_15_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_15_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_3_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_15_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_15_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_15_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_28_iswt1_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_15_a_core(nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_15_inst_ccs_lp_piped_fp_add_23_8_0_cmp_15_a_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_15_b_core(nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_15_inst_ccs_lp_piped_fp_add_23_8_0_cmp_15_b_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_15_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_15_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_15_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_1_cse)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_16 ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_16_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_16_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_5_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_16_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_16_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_16_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_28_oswt_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_16_a_core(ccs_lp_piped_fp_mult_23_8_0_cmp_25_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_16_b_core(nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_16_inst_ccs_lp_piped_fp_add_23_8_0_cmp_16_b_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_16_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_16_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_16_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_3_cse)
    );
  ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_17 ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_17_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_add_23_8_0_cmp_17_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_5_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_17_bawt(ccs_lp_piped_fp_add_23_8_0_cmp_17_bawt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_17_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_28_oswt_cse),
      .ccs_lp_piped_fp_add_23_8_0_cmp_17_a_core(ccs_lp_piped_fp_mult_23_8_0_cmp_27_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_17_b_core(nl_ist_core_ccs_lp_piped_fp_add_23_8_0_cmp_17_inst_ccs_lp_piped_fp_add_23_8_0_cmp_17_b_core[31:0]),
      .ccs_lp_piped_fp_add_23_8_0_cmp_17_z_mxwt(ccs_lp_piped_fp_add_23_8_0_cmp_17_z_mxwt),
      .ccs_lp_piped_fp_add_23_8_0_cmp_17_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_3_cse)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_3_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_28_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_a_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_b_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_1_cse)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1 ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_oswt_unreg(and_96_rmff),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_a_core(ccs_lp_piped_fp_recip_23_8_0_cmp_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_b_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_1_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_1_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_1_iswt1_pff(and_90_rmff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2 ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_oswt_unreg(and_96_rmff),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_a_core(ccs_lp_piped_fp_recip_23_8_0_cmp_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_b_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_2_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_2_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_2_iswt1_pff(and_90_rmff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_3 ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_3_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_oswt_unreg(and_96_rmff),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_3_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_a_core(ccs_lp_piped_fp_recip_23_8_0_cmp_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_b_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_3_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_3_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1_pff(and_90_rmff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4 ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_oswt_unreg(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_4_oswt_unreg),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1(ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_a_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_4_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_4_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_b_core(ist_req_stream_crt_sva_20_265_234),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_4_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1_pff(and_79_rmff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5 ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_oswt_unreg(and_77_rmff),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_5_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_a_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_5_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_b_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_5_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_5_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_5_iswt1_pff(and_76_rmff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6 ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_6_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_oswt_unreg(and_77_rmff),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_6_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_a_core(c_z_d_sva_12),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_b_core(n_z_d_sva_10),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_6_iswt1_pff(and_76_rmff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_7 ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_7_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_oswt_unreg(and_77_rmff),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_7_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_a_core(c_y_d_sva_12),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_b_core(n_y_d_sva_10),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_7_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_7_iswt1_pff(and_76_rmff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8 ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_8_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_oswt_unreg(and_77_rmff),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_8_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_a_core(c_x_d_sva_12),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_b_core(n_x_d_sva_10),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_8_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1_pff(and_76_rmff)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_9 ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_9_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_9_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_9_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_17_oswt_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_a_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_9_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_9_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_b_core(ccs_lp_piped_fp_add_23_8_0_cmp_10_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_9_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_7_cse)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10 ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_9_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_10_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_17_oswt_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_a_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_10_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_10_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_b_core(ccs_lp_piped_fp_add_23_8_0_cmp_11_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_10_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_10_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_7_cse)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_11 ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_11_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_9_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_11_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_17_oswt_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_a_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_11_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_11_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_b_core(ccs_lp_piped_fp_add_23_8_0_cmp_12_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_11_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_11_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_7_cse)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12 ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_9_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_12_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_17_oswt_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_a_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_12_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_12_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_b_core(ccs_lp_piped_fp_add_23_8_0_cmp_10_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_12_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_7_cse)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_13 ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_13_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_9_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_13_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_17_oswt_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_a_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_13_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_13_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_b_core(ccs_lp_piped_fp_add_23_8_0_cmp_11_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_13_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_13_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_7_cse)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14 ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_9_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_14_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_17_oswt_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_a_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_14_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_14_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_b_core(ccs_lp_piped_fp_add_23_8_0_cmp_12_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_14_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_14_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_7_cse)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_15 ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_15_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_7_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_15_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_a_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_15_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_15_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_b_core(ccs_lp_piped_fp_add_23_8_0_cmp_16_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_15_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_5_cse)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16 ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_7_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_16_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_a_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_16_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_16_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_b_core(ccs_lp_piped_fp_add_23_8_0_cmp_17_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_16_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_16_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_5_cse)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_17 ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_17_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_7_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_17_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_a_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_17_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_17_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_b_core(ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_17_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_17_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_5_cse)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18 ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_5_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_18_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_28_oswt_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_a_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_18_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_18_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_b_core(ccs_lp_piped_fp_add_23_8_0_cmp_15_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_18_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_18_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_3_cse)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_19 ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_19_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_5_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_19_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_28_oswt_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_a_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_19_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_19_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_b_core(ccs_lp_piped_fp_add_23_8_0_cmp_14_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_19_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_19_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_3_cse)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20 ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_5_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_20_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_28_oswt_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_a_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_20_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_20_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_b_core(ccs_lp_piped_fp_add_23_8_0_cmp_13_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_20_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_20_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_3_cse)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_21 ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_21_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_5_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_21_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_28_oswt_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_a_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_21_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_21_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_b_core(ccs_lp_piped_fp_add_23_8_0_cmp_15_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_21_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_21_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_3_cse)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22 ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_5_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_22_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_28_oswt_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_a_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_22_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_22_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_b_core(ccs_lp_piped_fp_add_23_8_0_cmp_14_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_22_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_22_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_3_cse)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_23 ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_23_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_5_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_23_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_28_oswt_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_a_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_23_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_23_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_b_core(ccs_lp_piped_fp_add_23_8_0_cmp_13_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_23_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_23_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_3_cse)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_24 ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_24_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_24_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_3_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_24_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_24_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_24_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_28_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_24_a_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_24_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_24_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_24_b_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_24_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_24_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_24_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_24_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_24_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_1_cse)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_25 ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_25_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_25_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_3_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_25_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_25_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_25_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_28_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_25_a_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_25_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_25_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_25_b_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_25_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_25_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_25_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_25_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_25_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_1_cse)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_26 ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_26_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_26_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_3_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_26_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_26_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_26_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_28_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_26_a_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_26_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_26_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_26_b_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_26_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_26_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_26_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_26_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_26_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_1_cse)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_27 ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_27_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_27_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_3_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_27_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_27_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_27_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_28_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_27_a_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_27_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_27_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_27_b_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_27_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_27_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_27_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_27_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_27_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_1_cse)
    );
  ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_28 ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_28_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_28_oswt_unreg(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_3_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_28_bawt(ccs_lp_piped_fp_mult_23_8_0_cmp_28_bawt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_28_iswt1(reg_ccs_lp_piped_fp_mult_23_8_0_cmp_28_iswt1_cse),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_28_a_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_28_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_28_a_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_28_b_core(nl_ist_core_ccs_lp_piped_fp_mult_23_8_0_cmp_28_inst_ccs_lp_piped_fp_mult_23_8_0_cmp_28_b_core[31:0]),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_28_z_mxwt(ccs_lp_piped_fp_mult_23_8_0_cmp_28_z_mxwt),
      .ccs_lp_piped_fp_mult_23_8_0_cmp_28_iswt1_pff(lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_1_cse)
    );
  ist_core_staller ist_core_staller_inst (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .core_wten(core_wten),
      .ist_req_stream_rsci_wen_comp(ist_req_stream_rsci_wen_comp),
      .ist_resp_stream_rsci_wen_comp(ist_resp_stream_rsci_wen_comp),
      .core_flen_unreg(nl_ist_core_staller_inst_core_flen_unreg)
    );
  ist_core_core_fsm ist_core_core_fsm_inst (
      .clk(clk),
      .arst_n(arst_n),
      .core_wen(core_wen),
      .fsm_output(fsm_output)
    );
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_15_mux1h_rmff = MUX_s_1_2_2(ccs_lp_piped_fp_add_23_8_0_cmp_3_b_core_31,
      operator_1_false_1_xor_tmp, and_31_tmp);
  assign nand_245_cse = ~(land_1_lpi_1_dfm_1_st_2 & main_stage_v_16);
  assign or_925_cse = ist_resp_stream_rsci_bawt | (~ reg_ist_resp_stream_rsci_iswt0_cse);
  assign or_924_cse = (~(main_stage_v_20 & land_1_lpi_1_dfm_1_st_6)) | ccs_lp_piped_fp_add_23_8_0_cmp_1_bawt;
  assign or_922_cse = (~(main_stage_v_18 & land_1_lpi_1_dfm_1_st_4)) | ccs_lp_piped_fp_add_23_8_0_cmp_2_bawt;
  assign or_920_cse = (~(main_stage_v_14 & land_lpi_1_dfm_2)) | ccs_lp_piped_fp_add_23_8_0_cmp_3_bawt;
  assign and_850_nl = nand_245_cse & and_tmp_26;
  assign and_851_nl = ccs_lp_piped_fp_mult_23_8_0_cmp_8_bawt & ccs_lp_piped_fp_mult_23_8_0_cmp_7_bawt
      & ccs_lp_piped_fp_mult_23_8_0_cmp_6_bawt & ccs_lp_piped_fp_mult_23_8_0_cmp_5_bawt;
  assign mux_167_nl = MUX_s_1_2_2(and_850_nl, and_tmp_26, and_851_nl);
  assign and_838_cse = mux_167_nl & or_925_cse & or_924_cse & or_922_cse & or_920_cse
      & ccs_lp_piped_fp_add_23_8_0_cmp_4_bawt & ccs_lp_piped_fp_add_23_8_0_cmp_6_bawt
      & main_stage_v_12 & core_wen;
  assign lp_piped_fp_add_AC_RND_CONV_0_32_8_15_mux1h_1_rmff = MUX_s_1_2_2(ccs_lp_piped_fp_add_23_8_0_cmp_3_a_core_31,
      operator_1_false_xor_tmp, and_31_tmp);
  assign and_632_cse = core_wen & (~ or_dcpl_5);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_1_cse
      = and_55_tmp & (fsm_output[1]);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_3_cse
      = and_51_tmp & (fsm_output[1]);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_5_cse
      = and_47_tmp & (fsm_output[1]);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_7_cse
      = and_43_tmp & (fsm_output[1]);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_9_cse
      = and_39_tmp & (fsm_output[1]);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_11_cse
      = and_35_tmp & (fsm_output[1]);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_13_cse
      = and_31_tmp & (fsm_output[1]);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_21_cse
      = and_15_tmp & (fsm_output[1]);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_20_cse
      = and_17_tmp & (fsm_output[1]);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_19_cse
      = and_19_tmp & (fsm_output[1]);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_18_cse
      = and_21_tmp & (fsm_output[1]);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_17_cse
      = and_23_tmp & (fsm_output[1]);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_16_cse
      = and_25_tmp & (fsm_output[1]);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_15_cse
      = and_27_tmp & (fsm_output[1]);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_14_cse
      = and_29_tmp & (fsm_output[1]);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_12_cse
      = and_33_tmp & (fsm_output[1]);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_10_cse
      = and_37_tmp & (fsm_output[1]);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_8_cse
      = and_41_tmp & (fsm_output[1]);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_6_cse
      = and_45_tmp & (fsm_output[1]);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_4_cse
      = and_49_tmp & (fsm_output[1]);
  assign lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_2_cse
      = and_53_tmp & (fsm_output[1]);
  assign and_76_rmff = mux_151_cse & land_lpi_1_dfm_2 & and_27_tmp;
  assign and_77_rmff = and_23_tmp & land_1_lpi_1_dfm_1_st_2;
  assign or_620_cse = ccs_fp_cmp_23_8_0_1_out_8 | ccs_fp_cmp_23_8_0_1_out_6;
  assign and_79_rmff = or_620_cse & and_764_cse;
  assign and_90_rmff = and_dcpl_20 & ccs_lp_piped_fp_recip_23_8_0_cmp_bawt & if_land_lpi_1_dfm_1_st_2
      & land_1_lpi_1_dfm_1_10 & main_stage_v_24;
  assign and_96_rmff = and_dcpl_25 & or_925_cse & ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt
      & if_land_lpi_1_dfm_1_st_4 & land_1_lpi_1_dfm_1_12 & main_stage_v_26;
  assign and_211_rmff = (~((ccs_lp_piped_fp_add_23_8_0_cmp_6_z_mxwt[31]) ^ (det_d_sva_2[31])))
      & (~((ccs_lp_piped_fp_add_23_8_0_cmp_4_z_mxwt[31]) ^ (det_d_sva_2[31]))) &
      and_31_tmp & (fsm_output[1]);
  assign and_100_rmff = and_19_tmp & land_1_lpi_1_dfm_1_st_4;
  assign and_106_rmff = FP_GEQ_32_8_lor_lpi_1_dfm_2 & if_land_lpi_1_dfm_2 & ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt
      & and_tmp_10 & or_925_cse & land_1_lpi_1_dfm_1_st_8 & main_stage_v_22;
  assign det_d_and_cse = core_wen & (~((~ mux_131_cse) | and_dcpl_4));
  assign and_743_cse = main_stage_v_22 & land_1_lpi_1_dfm_1_st_8;
  assign mux_83_nl = MUX_s_1_2_2(not_tmp_7, and_tmp_1, or_564_cse);
  assign and_58_nl = FP_GEQ_32_8_lor_lpi_1_dfm_st & land_1_lpi_1_dfm_1_st_7 & main_stage_v_21
      & mux_83_nl;
  assign or_562_nl = and_743_cse | and_tmp_1;
  assign mux_79_nl = MUX_s_1_2_2((~ nand_tmp_2), or_562_nl, and_744_cse);
  assign mux_82_nl = MUX_s_1_2_2((~ nand_tmp_2), mux_79_nl, FP_GEQ_32_8_lor_lpi_1_dfm_st);
  assign mux_84_nl = MUX_s_1_2_2(and_58_nl, mux_82_nl, FP_GEQ_32_8_lor_lpi_1_dfm_2);
  assign det_d_and_12_cse = det_d_and_cse & mux_84_nl;
  assign or_570_nl = (FP_GEQ_32_8_lor_lpi_1_dfm_2 & (~ ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt)
      & main_stage_v_22 & land_1_lpi_1_dfm_1_st_8) | and_tmp_4;
  assign mux_86_nl = MUX_s_1_2_2(nor_tmp_15, and_tmp_4, and_751_cse);
  assign or_569_nl = (~(ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt | (~ main_stage_v_22)
      | (~ land_1_lpi_1_dfm_1_st_8))) | and_tmp_4;
  assign mux_85_nl = MUX_s_1_2_2(and_743_cse, or_569_nl, and_751_cse);
  assign mux_87_nl = MUX_s_1_2_2(mux_86_nl, mux_85_nl, FP_GEQ_32_8_lor_lpi_1_dfm_2);
  assign mux_88_nl = MUX_s_1_2_2(or_570_nl, mux_87_nl, and_740_cse);
  assign mux_90_nl = MUX_s_1_2_2(mux_tmp_14, mux_88_nl, or_925_cse);
  assign mux_91_nl = MUX_s_1_2_2(mux_tmp_14, mux_90_nl, nand_217_cse);
  assign if_and_cse = det_d_and_cse & mux_91_nl;
  assign mux_105_nl = MUX_s_1_2_2(not_tmp_7, and_tmp_1, or_561_cse);
  assign and_765_nl = main_stage_v_22 & (~ mux_105_nl);
  assign or_576_nl = main_stage_v_22 | and_tmp_1;
  assign mux_106_nl = MUX_s_1_2_2(and_765_nl, or_576_nl, main_stage_v_21);
  assign FP_GEQ_32_8_oelse_and_cse = det_d_and_cse & mux_106_nl;
  assign and_642_cse = core_wen & (~ or_dcpl_20);
  assign and_767_nl = main_stage_v_24 & land_1_lpi_1_dfm_1_10 & if_land_lpi_1_dfm_1_st_2
      & (~(ccs_lp_piped_fp_recip_23_8_0_cmp_bawt & mux_tmp));
  assign or_578_nl = (main_stage_v_24 & land_1_lpi_1_dfm_1_10 & if_land_lpi_1_dfm_1_st_2)
      | mux_tmp;
  assign mux_107_nl = MUX_s_1_2_2(and_767_nl, or_578_nl, and_763_cse);
  assign and_799_cse = and_642_cse & mux_107_nl;
  assign if_aelse_and_2_cse = core_wen & (~ or_dcpl_30);
  assign mux_108_nl = MUX_s_1_2_2(or_925_cse, and_tmp, and_761_cse);
  assign and_771_nl = main_stage_v_26 & (~ mux_108_nl);
  assign or_579_nl = main_stage_v_26 | (~ reg_ist_resp_stream_rsci_iswt0_cse) | ist_resp_stream_rsci_bawt;
  assign mux_109_nl = MUX_s_1_2_2(and_771_nl, or_579_nl, main_stage_v_25);
  assign if_aelse_and_10_cse = if_aelse_and_2_cse & mux_109_nl;
  assign and_801_cse = core_wen & and_17_tmp & land_1_lpi_1_dfm_1_st_5;
  assign aelse_1_and_4_cse = core_wen & (~((~ and_17_tmp) | (fsm_output[0])));
  assign if_and_7_cse = core_wen & and_21_tmp & land_1_lpi_1_dfm_1_st_3;
  assign aelse_1_and_5_cse = core_wen & (~((~ and_21_tmp) | (fsm_output[0])));
  assign aelse_1_and_6_cse = core_wen & (~((~ and_25_tmp) | (fsm_output[0])));
  assign and_802_cse = core_wen & and_29_tmp & land_lpi_1_dfm_1;
  assign FP_LEQ_32_8_arelb_and_cse = core_wen & land_lpi_1_dfm_2 & and_27_tmp;
  assign aelse_and_cse = core_wen & (~((~ and_29_tmp) | (fsm_output[0])));
  assign det_d_and_3_cse = core_wen & (~((~ and_33_tmp) | (fsm_output[0])));
  assign and_660_cse = core_wen & (~((~ and_37_tmp) | (fsm_output[0])));
  assign and_664_cse = core_wen & (~((~ and_41_tmp) | (fsm_output[0])));
  assign and_667_cse = core_wen & (~((~ and_45_tmp) | (fsm_output[0])));
  assign and_670_cse = core_wen & (~((~ and_49_tmp) | (fsm_output[0])));
  assign and_673_cse = core_wen & (~((~ and_53_tmp) | (fsm_output[0])));
  assign det_d_and_4_cse = core_wen & and_15_tmp;
  assign mux_121_nl = MUX_s_1_2_2(not_tmp_23, or_tmp_34, and_751_cse);
  assign mux_122_nl = MUX_s_1_2_2(or_tmp_34, mux_121_nl, and_740_cse);
  assign mux_123_nl = MUX_s_1_2_2(not_tmp_23, mux_122_nl, or_925_cse);
  assign mux_124_nl = MUX_s_1_2_2(not_tmp_23, mux_123_nl, nand_217_cse);
  assign mux_125_nl = MUX_s_1_2_2((~ mux_124_nl), and_776_cse, and_15_tmp);
  assign det_d_and_15_cse = det_d_and_4_cse & mux_125_nl;
  assign mux_126_nl = MUX_s_1_2_2((~ FP_GEQ_32_8_lor_lpi_1_dfm_st), or_tmp_40, and_751_cse);
  assign mux_127_nl = MUX_s_1_2_2(or_tmp_40, mux_126_nl, and_740_cse);
  assign mux_128_nl = MUX_s_1_2_2(FP_GEQ_32_8_lor_lpi_1_dfm_st, (~ mux_127_nl), or_925_cse);
  assign mux_129_nl = MUX_s_1_2_2(FP_GEQ_32_8_lor_lpi_1_dfm_st, mux_128_nl, nand_217_cse);
  assign and_780_nl = main_stage_v_21 & land_1_lpi_1_dfm_1_st_7 & mux_129_nl;
  assign mux_130_nl = MUX_s_1_2_2(and_780_nl, and_776_cse, and_15_tmp);
  assign if_ttt_d_and_2_cse = det_d_and_4_cse & mux_130_nl;
  assign or_604_nl = and_763_cse | and_tmp_1;
  assign and_787_nl = if_land_lpi_1_dfm_2 & ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt
      & land_1_lpi_1_dfm_1_st_8;
  assign mux_166_nl = MUX_s_1_2_2(not_tmp_34, or_604_nl, and_787_nl);
  assign mux_136_nl = MUX_s_1_2_2(not_tmp_34, mux_166_nl, main_stage_v_22);
  assign mux_138_nl = MUX_s_1_2_2(not_tmp_34, mux_136_nl, FP_GEQ_32_8_lor_lpi_1_dfm_2);
  assign and_803_cse = and_642_cse & mux_138_nl;
  assign aelse_1_and_25_cse = and_642_cse & mux_tmp_66;
  assign or_608_nl = main_stage_v_25 | mux_tmp;
  assign mux_142_nl = MUX_s_1_2_2(not_tmp_39, or_608_nl, or_607_cse);
  assign mux_143_nl = MUX_s_1_2_2(not_tmp_39, mux_142_nl, main_stage_v_24);
  assign aelse_1_and_26_cse = if_aelse_and_2_cse & mux_143_nl;
  assign and_805_cse = core_wen & and_31_tmp & nor_105_cse;
  assign nor_105_cse = ~(operator_1_false_1_xor_tmp | operator_1_false_xor_tmp);
  assign and_806_cse = core_wen & and_19_tmp & land_1_lpi_1_dfm_1_st_4;
  assign and_679_cse = core_wen & (~((~ and_47_tmp) | (fsm_output[0])));
  assign and_680_cse = core_wen & (~((~ and_51_tmp) | (fsm_output[0])));
  assign and_681_cse = core_wen & (~((~ and_55_tmp) | (fsm_output[0])));
  assign and_682_cse = core_wen & (~((~ and_43_tmp) | (fsm_output[0])));
  assign det_d_and_7_cse = core_wen & (~((~ and_35_tmp) | (fsm_output[0])));
  assign and_683_cse = core_wen & (~((~ and_39_tmp) | (fsm_output[0])));
  assign aelse_and_2_cse = core_wen & (~((~ and_31_tmp) | (fsm_output[0])));
  assign if_and_10_cse = core_wen & and_23_tmp & land_1_lpi_1_dfm_1_st_2;
  assign aelse_1_and_11_cse = core_wen & (~((~ and_19_tmp) | (fsm_output[0])));
  assign aelse_1_and_12_cse = core_wen & (~((~ and_23_tmp) | (fsm_output[0])));
  assign aelse_1_and_13_cse = core_wen & (~((~ and_27_tmp) | (fsm_output[0])));
  assign FP_LEQ_32_8_FP_LEQ_32_8_or_cse = ccs_fp_cmp_23_8_0_out_7 | ccs_fp_cmp_23_8_0_out_6;
  assign and_791_nl = main_stage_v_24 & (~(or_607_cse & mux_tmp));
  assign or_610_nl = main_stage_v_24 | mux_tmp;
  assign mux_148_nl = MUX_s_1_2_2(and_791_nl, or_610_nl, main_stage_v_23);
  assign aelse_1_and_28_cse = and_642_cse & mux_148_nl;
  assign and_815_cse = core_wen & and_25_tmp & land_1_lpi_1_dfm_1_st_1;
  assign and_816_cse = core_wen & and_27_tmp & land_lpi_1_dfm_2 & mux_151_cse;
  assign operator_1_false_1_xor_tmp = (ccs_lp_piped_fp_add_23_8_0_cmp_4_z_mxwt[31])
      ^ (det_d_sva_2[31]);
  assign operator_1_false_xor_tmp = (ccs_lp_piped_fp_add_23_8_0_cmp_6_z_mxwt[31])
      ^ (det_d_sva_2[31]);
  assign nor_58_nl = ~(land_lpi_1_dfm_2 | (~(FP_LEQ_32_8_arelb_1_sva | fp_arelb_32_8_return_0_sva)));
  assign or_581_nl = land_lpi_1_dfm_2 | FP_LEQ_32_8_arelb_1_sva | fp_arelb_32_8_return_0_sva;
  assign mux_151_cse = MUX_s_1_2_2(nor_58_nl, or_581_nl, FP_LEQ_32_8_FP_LEQ_32_8_or_cse);
  assign and_55_tmp = ist_req_stream_rsci_bawt & or_369_cse_1 & or_370_cse_1 & or_371_cse_1
      & or_372_cse_1 & or_373_cse_1 & or_374_cse_1 & or_375_cse_1 & or_376_cse_1
      & or_377_cse_1 & or_289_cse_1 & or_290_cse_1 & or_291_cse_1 & or_292_cse_1
      & or_293_cse_1 & or_294_cse_1 & or_295_cse_1 & or_296_cse_1 & or_297_cse_1
      & or_227_cse_1 & or_228_cse_1 & or_229_cse_1 & or_230_cse_1 & or_231_cse_1
      & or_232_cse_1 & or_177_cse_1 & or_178_cse_1 & or_179_cse_1 & or_180_cse_1
      & or_181_cse_1 & or_182_cse_1 & or_183_cse_1 & or_141_cse_1 & or_142_cse_1
      & or_143_cse_1 & or_111_cse_1 & or_112_cse_1 & or_920_cse & or_61_cse_1 & or_62_cse_1
      & or_63_cse_1 & or_64_cse_1 & or_922_cse & or_924_cse & or_523_cse_1 & or_519_cse_1
      & or_1_cse_1 & or_2_cse_1 & or_3_cse_1 & or_925_cse;
  assign and_53_tmp = main_stage_v_1 & (~(main_stage_v_2 & (~ and_51_tmp))) & or_289_cse_1
      & or_290_cse_1 & or_291_cse_1 & or_292_cse_1 & or_293_cse_1 & or_294_cse_1
      & or_295_cse_1 & or_296_cse_1 & or_297_cse_1 & or_227_cse_1 & or_228_cse_1
      & or_229_cse_1 & or_230_cse_1 & or_231_cse_1 & or_232_cse_1 & or_177_cse_1
      & or_178_cse_1 & or_179_cse_1 & or_180_cse_1 & or_181_cse_1 & or_182_cse_1
      & or_183_cse_1 & or_141_cse_1 & or_142_cse_1 & or_143_cse_1 & or_111_cse_1
      & or_112_cse_1 & or_920_cse & or_61_cse_1 & or_62_cse_1 & or_63_cse_1 & or_64_cse_1
      & or_922_cse & or_924_cse & or_523_cse_1 & or_519_cse_1 & or_1_cse_1 & or_2_cse_1
      & or_3_cse_1 & or_925_cse;
  assign and_51_tmp = main_stage_v_2 & or_369_cse_1 & or_370_cse_1 & or_371_cse_1
      & or_372_cse_1 & or_373_cse_1 & or_374_cse_1 & or_375_cse_1 & or_376_cse_1
      & or_377_cse_1 & or_289_cse_1 & or_290_cse_1 & or_291_cse_1 & or_292_cse_1
      & or_293_cse_1 & or_294_cse_1 & or_295_cse_1 & or_296_cse_1 & or_297_cse_1
      & or_227_cse_1 & or_228_cse_1 & or_229_cse_1 & or_230_cse_1 & or_231_cse_1
      & or_232_cse_1 & or_177_cse_1 & or_178_cse_1 & or_179_cse_1 & or_180_cse_1
      & or_181_cse_1 & or_182_cse_1 & or_183_cse_1 & or_141_cse_1 & or_142_cse_1
      & or_143_cse_1 & or_111_cse_1 & or_112_cse_1 & or_920_cse & or_61_cse_1 & or_62_cse_1
      & or_63_cse_1 & or_64_cse_1 & or_922_cse & or_924_cse & or_523_cse_1 & or_519_cse_1
      & or_1_cse_1 & or_2_cse_1 & or_3_cse_1 & or_925_cse;
  assign and_49_tmp = main_stage_v_3 & (~(main_stage_v_4 & (~ and_47_tmp))) & or_227_cse_1
      & or_228_cse_1 & or_229_cse_1 & or_230_cse_1 & or_231_cse_1 & or_232_cse_1
      & or_177_cse_1 & or_178_cse_1 & or_179_cse_1 & or_180_cse_1 & or_181_cse_1
      & or_182_cse_1 & or_183_cse_1 & or_141_cse_1 & or_142_cse_1 & or_143_cse_1
      & or_111_cse_1 & or_112_cse_1 & or_920_cse & or_61_cse_1 & or_62_cse_1 & or_63_cse_1
      & or_64_cse_1 & or_922_cse & or_924_cse & or_523_cse_1 & or_519_cse_1 & or_1_cse_1
      & or_2_cse_1 & or_3_cse_1 & or_925_cse;
  assign and_47_tmp = main_stage_v_4 & or_289_cse_1 & or_290_cse_1 & or_291_cse_1
      & or_292_cse_1 & or_293_cse_1 & or_294_cse_1 & or_295_cse_1 & or_296_cse_1
      & or_297_cse_1 & or_227_cse_1 & or_228_cse_1 & or_229_cse_1 & or_230_cse_1
      & or_231_cse_1 & or_232_cse_1 & or_177_cse_1 & or_178_cse_1 & or_179_cse_1
      & or_180_cse_1 & or_181_cse_1 & or_182_cse_1 & or_183_cse_1 & or_141_cse_1
      & or_142_cse_1 & or_143_cse_1 & or_111_cse_1 & or_112_cse_1 & or_920_cse &
      or_61_cse_1 & or_62_cse_1 & or_63_cse_1 & or_64_cse_1 & or_922_cse & or_924_cse
      & or_523_cse_1 & or_519_cse_1 & or_1_cse_1 & or_2_cse_1 & or_3_cse_1 & or_925_cse;
  assign and_45_tmp = main_stage_v_5 & (~(main_stage_v_6 & (~ and_43_tmp))) & or_177_cse_1
      & or_178_cse_1 & or_179_cse_1 & or_180_cse_1 & or_181_cse_1 & or_182_cse_1
      & or_183_cse_1 & or_141_cse_1 & or_142_cse_1 & or_143_cse_1 & or_111_cse_1
      & or_112_cse_1 & or_920_cse & or_61_cse_1 & or_62_cse_1 & or_63_cse_1 & or_64_cse_1
      & or_922_cse & or_924_cse & or_523_cse_1 & or_519_cse_1 & or_1_cse_1 & or_2_cse_1
      & or_3_cse_1 & or_925_cse;
  assign and_43_tmp = main_stage_v_6 & or_227_cse_1 & or_228_cse_1 & or_229_cse_1
      & or_230_cse_1 & or_231_cse_1 & or_232_cse_1 & or_177_cse_1 & or_178_cse_1
      & or_179_cse_1 & or_180_cse_1 & or_181_cse_1 & or_182_cse_1 & or_183_cse_1
      & or_141_cse_1 & or_142_cse_1 & or_143_cse_1 & or_111_cse_1 & or_112_cse_1
      & or_920_cse & or_61_cse_1 & or_62_cse_1 & or_63_cse_1 & or_64_cse_1 & or_922_cse
      & or_924_cse & or_523_cse_1 & or_519_cse_1 & or_1_cse_1 & or_2_cse_1 & or_3_cse_1
      & or_925_cse;
  assign and_41_tmp = main_stage_v_7 & (~(main_stage_v_8 & (~ and_39_tmp))) & or_141_cse_1
      & or_142_cse_1 & or_143_cse_1 & or_111_cse_1 & or_112_cse_1 & or_920_cse &
      or_61_cse_1 & or_62_cse_1 & or_63_cse_1 & or_64_cse_1 & or_922_cse & or_924_cse
      & or_523_cse_1 & or_519_cse_1 & or_1_cse_1 & or_2_cse_1 & or_3_cse_1 & or_925_cse;
  assign and_39_tmp = main_stage_v_8 & or_177_cse_1 & or_178_cse_1 & or_179_cse_1
      & or_180_cse_1 & or_181_cse_1 & or_182_cse_1 & or_183_cse_1 & or_141_cse_1
      & or_142_cse_1 & or_143_cse_1 & or_111_cse_1 & or_112_cse_1 & or_920_cse &
      or_61_cse_1 & or_62_cse_1 & or_63_cse_1 & or_64_cse_1 & or_922_cse & or_924_cse
      & or_523_cse_1 & or_519_cse_1 & or_1_cse_1 & or_2_cse_1 & or_3_cse_1 & or_925_cse;
  assign and_37_tmp = main_stage_v_9 & (~(main_stage_v_10 & (~ and_35_tmp))) & or_111_cse_1
      & or_112_cse_1 & or_920_cse & or_61_cse_1 & or_62_cse_1 & or_63_cse_1 & or_64_cse_1
      & or_922_cse & or_924_cse & or_523_cse_1 & or_519_cse_1 & or_1_cse_1 & or_2_cse_1
      & or_3_cse_1 & or_925_cse;
  assign and_35_tmp = main_stage_v_10 & or_141_cse_1 & or_142_cse_1 & or_143_cse_1
      & or_111_cse_1 & or_112_cse_1 & or_920_cse & or_61_cse_1 & or_62_cse_1 & or_63_cse_1
      & or_64_cse_1 & or_922_cse & or_924_cse & or_523_cse_1 & or_519_cse_1 & or_1_cse_1
      & or_2_cse_1 & or_3_cse_1 & or_925_cse;
  assign and_33_tmp = main_stage_v_11 & or_111_cse_1 & or_112_cse_1 & or_920_cse
      & or_61_cse_1 & or_62_cse_1 & or_63_cse_1 & or_64_cse_1 & or_922_cse & or_924_cse
      & or_523_cse_1 & or_519_cse_1 & or_1_cse_1 & or_2_cse_1 & or_3_cse_1 & or_925_cse;
  assign and_31_tmp = main_stage_v_12 & or_111_cse_1 & or_112_cse_1 & or_920_cse
      & or_61_cse_1 & or_62_cse_1 & or_63_cse_1 & or_64_cse_1 & or_922_cse & or_924_cse
      & or_523_cse_1 & or_519_cse_1 & or_1_cse_1 & or_2_cse_1 & or_3_cse_1 & or_925_cse;
  assign and_29_tmp = main_stage_v_13 & or_920_cse & or_61_cse_1 & or_62_cse_1 &
      or_63_cse_1 & or_64_cse_1 & or_922_cse & or_924_cse & or_523_cse_1 & or_519_cse_1
      & or_1_cse_1 & or_2_cse_1 & or_3_cse_1 & or_925_cse;
  assign and_27_tmp = main_stage_v_14 & or_920_cse & or_61_cse_1 & or_62_cse_1 &
      or_63_cse_1 & or_64_cse_1 & or_922_cse & or_924_cse & or_523_cse_1 & or_519_cse_1
      & or_1_cse_1 & or_2_cse_1 & or_3_cse_1 & or_925_cse;
  assign and_25_tmp = main_stage_v_15 & or_61_cse_1 & or_62_cse_1 & or_63_cse_1 &
      or_64_cse_1 & or_922_cse & or_924_cse & or_523_cse_1 & or_519_cse_1 & or_1_cse_1
      & or_2_cse_1 & or_3_cse_1 & or_925_cse;
  assign and_23_tmp = main_stage_v_16 & or_61_cse_1 & or_62_cse_1 & or_63_cse_1 &
      or_64_cse_1 & or_922_cse & or_924_cse & or_523_cse_1 & or_519_cse_1 & or_1_cse_1
      & or_2_cse_1 & or_3_cse_1 & or_925_cse;
  assign and_21_tmp = main_stage_v_17 & or_922_cse & or_924_cse & or_523_cse_1 &
      or_519_cse_1 & or_1_cse_1 & or_2_cse_1 & or_3_cse_1 & or_925_cse;
  assign and_19_tmp = main_stage_v_18 & or_922_cse & or_924_cse & or_523_cse_1 &
      or_519_cse_1 & or_1_cse_1 & or_2_cse_1 & or_3_cse_1 & or_925_cse;
  assign and_17_tmp = main_stage_v_19 & or_924_cse & or_523_cse_1 & or_519_cse_1
      & or_1_cse_1 & or_2_cse_1 & or_3_cse_1 & or_925_cse;
  assign and_15_tmp = main_stage_v_20 & or_924_cse & or_523_cse_1 & or_519_cse_1
      & or_1_cse_1 & or_2_cse_1 & or_3_cse_1 & or_925_cse;
  assign operator_1_false_return_2_sva_mx0w0 = (ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt[31])
      ^ (det_d_sva_10[31]);
  assign if_land_lpi_1_dfm_1_mx0w0 = if_land_lpi_1_dfm_2 & FP_GEQ_32_8_lor_lpi_1_dfm_2;
  assign if_land_lpi_1_dfm_2 = ccs_fp_cmp_23_8_0_2_out_7 | ccs_fp_cmp_23_8_0_2_out_6;
  assign or_369_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_bawt | (~ main_stage_v_2);
  assign or_370_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_28_bawt | (~ main_stage_v_2);
  assign or_371_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_27_bawt | (~ main_stage_v_2);
  assign or_372_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_26_bawt | (~ main_stage_v_2);
  assign or_373_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_25_bawt | (~ main_stage_v_2);
  assign or_374_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_24_bawt | (~ main_stage_v_2);
  assign or_375_cse_1 = ccs_lp_piped_fp_add_23_8_0_cmp_15_bawt | (~ main_stage_v_2);
  assign or_376_cse_1 = ccs_lp_piped_fp_add_23_8_0_cmp_14_bawt | (~ main_stage_v_2);
  assign or_377_cse_1 = ccs_lp_piped_fp_add_23_8_0_cmp_13_bawt | (~ main_stage_v_2);
  assign or_289_cse_1 = ccs_lp_piped_fp_add_23_8_0_cmp_bawt | (~ main_stage_v_4);
  assign or_290_cse_1 = ccs_lp_piped_fp_add_23_8_0_cmp_17_bawt | (~ main_stage_v_4);
  assign or_291_cse_1 = ccs_lp_piped_fp_add_23_8_0_cmp_16_bawt | (~ main_stage_v_4);
  assign or_292_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_23_bawt | (~ main_stage_v_4);
  assign or_293_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_22_bawt | (~ main_stage_v_4);
  assign or_294_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_21_bawt | (~ main_stage_v_4);
  assign or_295_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_20_bawt | (~ main_stage_v_4);
  assign or_296_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_19_bawt | (~ main_stage_v_4);
  assign or_297_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_18_bawt | (~ main_stage_v_4);
  assign or_227_cse_1 = ccs_lp_piped_fp_add_23_8_0_cmp_12_bawt | (~ main_stage_v_6);
  assign or_228_cse_1 = ccs_lp_piped_fp_add_23_8_0_cmp_11_bawt | (~ main_stage_v_6);
  assign or_229_cse_1 = ccs_lp_piped_fp_add_23_8_0_cmp_10_bawt | (~ main_stage_v_6);
  assign or_230_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_17_bawt | (~ main_stage_v_6);
  assign or_231_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_16_bawt | (~ main_stage_v_6);
  assign or_232_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_15_bawt | (~ main_stage_v_6);
  assign or_177_cse_1 = ccs_lp_piped_fp_add_23_8_0_cmp_9_bawt | (~ main_stage_v_8);
  assign or_178_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_14_bawt | (~ main_stage_v_8);
  assign or_179_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_13_bawt | (~ main_stage_v_8);
  assign or_180_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_12_bawt | (~ main_stage_v_8);
  assign or_181_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_11_bawt | (~ main_stage_v_8);
  assign or_182_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_10_bawt | (~ main_stage_v_8);
  assign or_183_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_9_bawt | (~ main_stage_v_8);
  assign or_141_cse_1 = ccs_lp_piped_fp_add_23_8_0_cmp_8_bawt | (~ main_stage_v_10);
  assign or_142_cse_1 = ccs_lp_piped_fp_add_23_8_0_cmp_7_bawt | (~ main_stage_v_10);
  assign or_143_cse_1 = ccs_lp_piped_fp_add_23_8_0_cmp_5_bawt | (~ main_stage_v_10);
  assign or_111_cse_1 = ccs_lp_piped_fp_add_23_8_0_cmp_6_bawt | (~ main_stage_v_12);
  assign or_112_cse_1 = ccs_lp_piped_fp_add_23_8_0_cmp_4_bawt | (~ main_stage_v_12);
  assign or_61_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_8_bawt | nand_245_cse;
  assign or_62_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_7_bawt | nand_245_cse;
  assign or_63_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_6_bawt | nand_245_cse;
  assign or_64_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_5_bawt | nand_245_cse;
  assign or_523_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt | (~(FP_GEQ_32_8_lor_lpi_1_dfm_2
      & land_1_lpi_1_dfm_1_st_8 & main_stage_v_22));
  assign or_519_cse_1 = ccs_lp_piped_fp_recip_23_8_0_cmp_bawt | (~(if_land_lpi_1_dfm_1_st_2
      & land_1_lpi_1_dfm_1_10 & main_stage_v_24));
  assign or_1_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_3_bawt | nand_5_cse_1;
  assign or_2_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt | nand_5_cse_1;
  assign or_3_cse_1 = ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt | nand_5_cse_1;
  assign nand_5_cse_1 = ~(if_land_lpi_1_dfm_1_st_4 & land_1_lpi_1_dfm_1_12 & main_stage_v_26);
  assign and_tmp = ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt & ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt
      & ccs_lp_piped_fp_mult_23_8_0_cmp_3_bawt & or_925_cse;
  assign and_740_cse = main_stage_v_26 & land_1_lpi_1_dfm_1_12 & if_land_lpi_1_dfm_1_st_4;
  assign mux_tmp = MUX_s_1_2_2(or_925_cse, and_tmp, and_740_cse);
  assign nand_217_cse = ~(main_stage_v_24 & land_1_lpi_1_dfm_1_10 & if_land_lpi_1_dfm_1_st_2
      & (~ ccs_lp_piped_fp_recip_23_8_0_cmp_bawt));
  assign and_tmp_1 = nand_217_cse & mux_tmp;
  assign or_561_cse = (~ FP_GEQ_32_8_lor_lpi_1_dfm_2) | ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt;
  assign and_797_nl = land_1_lpi_1_dfm_1_st_8 & (~ and_tmp_1);
  assign mux_78_nl = MUX_s_1_2_2(land_1_lpi_1_dfm_1_st_8, and_797_nl, ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt);
  assign nand_tmp_2 = ~(main_stage_v_22 & FP_GEQ_32_8_lor_lpi_1_dfm_2 & mux_78_nl);
  assign not_tmp_7 = ~(land_1_lpi_1_dfm_1_st_8 | (~ and_tmp_1));
  assign or_564_cse = (~ main_stage_v_22) | (~ FP_GEQ_32_8_lor_lpi_1_dfm_2) | ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt;
  assign and_744_cse = land_1_lpi_1_dfm_1_st_7 & main_stage_v_21;
  assign and_tmp_4 = main_stage_v_21 & land_1_lpi_1_dfm_1_st_7 & FP_GEQ_32_8_lor_lpi_1_dfm_st;
  assign nor_tmp_15 = FP_GEQ_32_8_lor_lpi_1_dfm_2 & main_stage_v_22 & land_1_lpi_1_dfm_1_st_8;
  assign mux_tmp_14 = MUX_s_1_2_2(nor_tmp_15, and_743_cse, FP_GEQ_32_8_lor_lpi_1_dfm_2);
  assign and_751_cse = ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt & ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt
      & ccs_lp_piped_fp_mult_23_8_0_cmp_3_bawt;
  assign or_tmp_15 = and_743_cse | (~ reg_ist_resp_stream_rsci_iswt0_cse) | ist_resp_stream_rsci_bawt;
  assign nand_tmp_3 = ~(main_stage_v_22 & land_1_lpi_1_dfm_1_st_8 & (~(or_561_cse
      & or_925_cse)));
  assign mux_94_nl = MUX_s_1_2_2(and_743_cse, (~ nand_tmp_3), and_751_cse);
  assign mux_92_nl = MUX_s_1_2_2((~ nand_tmp_3), or_tmp_15, land_1_lpi_1_dfm_1_st_7);
  assign mux_93_nl = MUX_s_1_2_2(and_743_cse, mux_92_nl, and_751_cse);
  assign mux_tmp_20 = MUX_s_1_2_2(mux_94_nl, mux_93_nl, main_stage_v_21);
  assign mux_tmp_21 = MUX_s_1_2_2((~ nand_tmp_3), or_tmp_15, and_744_cse);
  assign mux_tmp_22 = MUX_s_1_2_2(mux_tmp_21, mux_tmp_20, and_740_cse);
  assign and_763_cse = main_stage_v_23 & if_land_lpi_1_dfm_1_st_1 & land_1_lpi_1_dfm_1_st_9;
  assign and_761_cse = land_1_lpi_1_dfm_1_12 & if_land_lpi_1_dfm_1_st_4;
  assign and_764_cse = land_1_lpi_1_dfm_1_st_6 & and_15_tmp;
  assign not_tmp_23 = ~(main_stage_v_21 & land_1_lpi_1_dfm_1_st_7 & FP_GEQ_32_8_lor_lpi_1_dfm_st);
  assign nand_223_cse = ~(main_stage_v_22 & land_1_lpi_1_dfm_1_st_8 & FP_GEQ_32_8_lor_lpi_1_dfm_2
      & (~ ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt));
  assign or_tmp_34 = nand_223_cse | not_tmp_23;
  assign and_776_cse = or_620_cse & land_1_lpi_1_dfm_1_st_6;
  assign or_tmp_40 = nand_223_cse | (~ FP_GEQ_32_8_lor_lpi_1_dfm_st);
  assign nand_228_cse = ~(ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt & ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt
      & ccs_lp_piped_fp_mult_23_8_0_cmp_3_bawt);
  assign nand_206_cse = ~(main_stage_v_26 & land_1_lpi_1_dfm_1_12 & if_land_lpi_1_dfm_1_st_4
      & nand_228_cse);
  assign and_tmp_10 = nand_217_cse & nand_206_cse;
  assign nor_56_nl = ~(land_1_lpi_1_dfm_1_st_8 | (~ and_tmp_10));
  assign mux_131_cse = MUX_s_1_2_2(nor_56_nl, and_tmp_10, or_564_cse);
  assign not_tmp_34 = land_1_lpi_1_dfm_1_st_9 & if_land_lpi_1_dfm_1_st_1 & main_stage_v_23
      & (~ and_tmp_1);
  assign or_tmp_47 = main_stage_v_23 | and_tmp_1;
  assign nand_tmp_11 = ~(main_stage_v_23 & (~ and_tmp_1));
  assign mux_139_nl = MUX_s_1_2_2(or_tmp_47, (~ nand_tmp_11), land_1_lpi_1_dfm_1_st_8);
  assign mux_140_nl = MUX_s_1_2_2(mux_139_nl, or_tmp_47, or_561_cse);
  assign mux_tmp_66 = MUX_s_1_2_2((~ nand_tmp_11), mux_140_nl, main_stage_v_22);
  assign not_tmp_39 = main_stage_v_25 & (~ mux_tmp);
  assign or_607_cse = (~ land_1_lpi_1_dfm_1_10) | (~ if_land_lpi_1_dfm_1_st_2) |
      ccs_lp_piped_fp_recip_23_8_0_cmp_bawt;
  assign and_dcpl_4 = (~ ist_resp_stream_rsci_bawt) & reg_ist_resp_stream_rsci_iswt0_cse;
  assign and_dcpl_6 = nand_228_cse & and_761_cse;
  assign or_dcpl_5 = and_dcpl_6 | and_dcpl_4 | (~ main_stage_v_26);
  assign and_dcpl_15 = and_tmp_10 & or_925_cse;
  assign and_dcpl_20 = nand_206_cse & or_925_cse;
  assign and_dcpl_25 = ccs_lp_piped_fp_mult_23_8_0_cmp_3_bawt & ccs_lp_piped_fp_mult_23_8_0_cmp_2_bawt;
  assign and_dcpl_37 = ((and_dcpl_25 & ccs_lp_piped_fp_mult_23_8_0_cmp_1_bawt) |
      (~(if_land_lpi_1_dfm_1_st_4 & land_1_lpi_1_dfm_1_12))) & or_925_cse;
  assign and_dcpl_39 = ist_resp_stream_rsci_bawt & reg_ist_resp_stream_rsci_iswt0_cse;
  assign and_dcpl_40 = (and_dcpl_6 | (~ main_stage_v_26)) & and_dcpl_39;
  assign and_dcpl_42 = mux_131_cse & or_925_cse;
  assign and_dcpl_47 = and_dcpl_15 & ((~ land_1_lpi_1_dfm_1_st_8) | ccs_lp_piped_fp_mult_23_8_0_cmp_4_bawt
      | (~ FP_GEQ_32_8_lor_lpi_1_dfm_2));
  assign or_dcpl_20 = (~ and_tmp_10) | and_dcpl_4;
  assign or_dcpl_25 = (~ and_tmp_10) | and_dcpl_4 | (~ main_stage_v_23);
  assign and_dcpl_56 = and_dcpl_20 & or_607_cse;
  assign and_dcpl_61 = nand_228_cse & and_761_cse & main_stage_v_26;
  assign or_dcpl_30 = and_dcpl_61 | and_dcpl_4;
  assign or_dcpl_34 = and_dcpl_61 | and_dcpl_4 | (~ main_stage_v_25);
  assign and_dcpl_110 = and_dcpl_15 & (~ land_1_lpi_1_dfm_1_st_8);
  assign main_stage_v_21_mx0c1 = and_dcpl_42 & main_stage_v_21 & (~ and_15_tmp);
  assign main_stage_v_22_mx0c1 = and_dcpl_47 & main_stage_v_22 & (~ main_stage_v_21);
  assign nor_59_nl = ~(or_561_cse | (~(land_1_lpi_1_dfm_1_st_8 & and_tmp_10)));
  assign mux_160_nl = MUX_s_1_2_2(and_tmp_10, nor_59_nl, main_stage_v_22);
  assign main_stage_v_23_mx0c1 = mux_160_nl & or_925_cse & main_stage_v_23;
  assign main_stage_v_24_mx0c1 = and_dcpl_56 & main_stage_v_24 & (~ main_stage_v_23);
  assign or_656_nl = or_607_cse | and_dcpl_61;
  assign mux_163_nl = MUX_s_1_2_2(and_dcpl_61, or_656_nl, main_stage_v_24);
  assign main_stage_v_25_mx0c1 = (~ mux_163_nl) & or_925_cse & main_stage_v_25;
  assign main_stage_v_26_mx0c1 = and_dcpl_37 & main_stage_v_26 & (~ main_stage_v_25);
  assign main_stage_v_20_mx0c1 = and_15_tmp & (~ and_17_tmp) & (fsm_output[1]);
  assign main_stage_v_19_mx0c1 = (~ and_19_tmp) & and_17_tmp & (fsm_output[1]);
  assign main_stage_v_18_mx0c1 = and_19_tmp & (~ and_21_tmp) & (fsm_output[1]);
  assign main_stage_v_17_mx0c1 = (~ and_23_tmp) & and_21_tmp & (fsm_output[1]);
  assign main_stage_v_16_mx0c1 = and_23_tmp & (~ and_25_tmp) & (fsm_output[1]);
  assign main_stage_v_15_mx0c1 = (~ and_27_tmp) & and_25_tmp & (fsm_output[1]);
  assign main_stage_v_14_mx0c1 = and_27_tmp & (~ and_29_tmp) & (fsm_output[1]);
  assign main_stage_v_13_mx0c1 = (~ and_31_tmp) & and_29_tmp & (fsm_output[1]);
  assign main_stage_v_12_mx0c1 = and_31_tmp & (~ and_33_tmp) & (fsm_output[1]);
  assign main_stage_v_11_mx0c1 = (~ and_35_tmp) & and_33_tmp & (fsm_output[1]);
  assign main_stage_v_10_mx0c1 = (~ and_37_tmp) & and_35_tmp & (fsm_output[1]);
  assign main_stage_v_9_mx0c1 = (~ and_39_tmp) & and_37_tmp & (fsm_output[1]);
  assign main_stage_v_8_mx0c1 = and_39_tmp & (~ and_41_tmp) & (fsm_output[1]);
  assign main_stage_v_7_mx0c1 = (~ and_43_tmp) & and_41_tmp & (fsm_output[1]);
  assign main_stage_v_6_mx0c1 = and_43_tmp & (~ and_45_tmp) & (fsm_output[1]);
  assign main_stage_v_5_mx0c1 = (~ and_47_tmp) & and_45_tmp & (fsm_output[1]);
  assign main_stage_v_4_mx0c1 = (~ and_49_tmp) & and_47_tmp & (fsm_output[1]);
  assign main_stage_v_3_mx0c1 = and_49_tmp & (~ and_51_tmp) & (fsm_output[1]);
  assign main_stage_v_2_mx0c1 = (~ and_53_tmp) & and_51_tmp & (fsm_output[1]);
  assign main_stage_v_1_mx0c1 = and_53_tmp & (~ and_55_tmp) & (fsm_output[1]);
  assign and_tmp_26 = nand_223_cse & nand_217_cse & (and_751_cse | nand_5_cse_1);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ist_req_stream_rsci_iswt0 <= 1'b0;
    end
    else if ( core_wen & (and_55_tmp | (fsm_output[0])) ) begin
      ist_req_stream_rsci_iswt0 <= 1'b1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_3_b_core_31 <= 1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_3_a_core_31 <= 1'b0;
    end
    else if ( and_838_cse ) begin
      ccs_lp_piped_fp_add_23_8_0_cmp_3_b_core_31 <= lp_piped_fp_add_AC_RND_CONV_0_32_8_15_mux1h_rmff;
      ccs_lp_piped_fp_add_23_8_0_cmp_3_a_core_31 <= lp_piped_fp_add_AC_RND_CONV_0_32_8_15_mux1h_1_rmff;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ist_resp_stream_rsci_idat_9_0 <= 10'b0000000000;
      ist_resp_stream_rsci_idat_10 <= 1'b0;
      ist_resp_stream_rsci_idat_42_11 <= 32'b00000000000000000000000000000000;
      ist_resp_stream_rsci_idat_74_43 <= 32'b00000000000000000000000000000000;
      ist_resp_stream_rsci_idat_106_75 <= 32'b00000000000000000000000000000000;
    end
    else if ( and_632_cse ) begin
      ist_resp_stream_rsci_idat_9_0 <= ist_req_stream_rid_slc_ist_req_stream_crt_9_0_itm_6;
      ist_resp_stream_rsci_idat_10 <= if_if_if_if_and_itm_4;
      ist_resp_stream_rsci_idat_42_11 <= ccs_lp_piped_fp_mult_23_8_0_cmp_3_z_mxwt
          & ({{31{if_land_lpi_1_dfm_1_st_4}}, if_land_lpi_1_dfm_1_st_4}) & ({{31{land_1_lpi_1_dfm_1_12}},
          land_1_lpi_1_dfm_1_12});
      ist_resp_stream_rsci_idat_74_43 <= ccs_lp_piped_fp_mult_23_8_0_cmp_2_z_mxwt
          & ({{31{if_land_lpi_1_dfm_1_st_4}}, if_land_lpi_1_dfm_1_st_4}) & ({{31{land_1_lpi_1_dfm_1_12}},
          land_1_lpi_1_dfm_1_12});
      ist_resp_stream_rsci_idat_106_75 <= ccs_lp_piped_fp_mult_23_8_0_cmp_1_z_mxwt
          & ({{31{if_land_lpi_1_dfm_1_st_4}}, if_land_lpi_1_dfm_1_st_4}) & ({{31{land_1_lpi_1_dfm_1_12}},
          land_1_lpi_1_dfm_1_12});
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_ccs_lp_piped_fp_mult_23_8_0_cmp_28_iswt1_cse <= 1'b0;
      reg_ccs_lp_piped_fp_mult_23_8_0_cmp_28_oswt_cse <= 1'b0;
      reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_cse <= 1'b0;
      reg_ccs_lp_piped_fp_mult_23_8_0_cmp_17_oswt_cse <= 1'b0;
      reg_ccs_lp_piped_fp_mult_23_8_0_cmp_14_oswt_cse <= 1'b0;
      reg_ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1_cse <= 1'b0;
      reg_ccs_lp_piped_fp_mult_23_8_0_cmp_8_oswt_cse <= 1'b0;
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1 <= 1'b0;
      reg_ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1_cse <= 1'b0;
      reg_ccs_lp_piped_fp_add_23_8_0_cmp_8_oswt_cse <= 1'b0;
      ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1 <= 1'b0;
      reg_ccs_lp_piped_fp_add_23_8_0_cmp_2_oswt_cse <= 1'b0;
      ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1 <= 1'b0;
    end
    else if ( core_wen ) begin
      reg_ccs_lp_piped_fp_mult_23_8_0_cmp_28_iswt1_cse <= lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_1_cse;
      reg_ccs_lp_piped_fp_mult_23_8_0_cmp_28_oswt_cse <= lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_3_cse;
      reg_ccs_lp_piped_fp_mult_23_8_0_cmp_23_oswt_cse <= lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_5_cse;
      reg_ccs_lp_piped_fp_mult_23_8_0_cmp_17_oswt_cse <= lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_7_cse;
      reg_ccs_lp_piped_fp_mult_23_8_0_cmp_14_oswt_cse <= lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_9_cse;
      reg_ccs_lp_piped_fp_mult_23_8_0_cmp_8_iswt1_cse <= and_76_rmff;
      reg_ccs_lp_piped_fp_mult_23_8_0_cmp_8_oswt_cse <= and_77_rmff;
      ccs_lp_piped_fp_mult_23_8_0_cmp_4_iswt1 <= and_79_rmff;
      reg_ccs_lp_piped_fp_mult_23_8_0_cmp_3_iswt1_cse <= and_90_rmff;
      reg_ccs_lp_piped_fp_add_23_8_0_cmp_8_oswt_cse <= lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_11_cse;
      ccs_lp_piped_fp_add_23_8_0_cmp_3_iswt1 <= and_211_rmff;
      reg_ccs_lp_piped_fp_add_23_8_0_cmp_2_oswt_cse <= and_100_rmff;
      ccs_lp_piped_fp_recip_23_8_0_cmp_iswt1 <= and_106_rmff;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_ist_resp_stream_rsci_iswt0_cse <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_37 & main_stage_v_26) | and_dcpl_40) ) begin
      reg_ist_resp_stream_rsci_iswt0_cse <= ~ and_dcpl_40;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_21 <= 1'b0;
    end
    else if ( core_wen & (lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_21_cse
        | main_stage_v_21_mx0c1) ) begin
      main_stage_v_21 <= ~ main_stage_v_21_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_22 <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_42 & main_stage_v_21) | main_stage_v_22_mx0c1)
        ) begin
      main_stage_v_22 <= ~ main_stage_v_22_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      det_d_sva_12_30_0 <= 31'b0000000000000000000000000000000;
      operator_1_false_return_sva_10 <= 1'b0;
      operator_1_false_return_1_sva_10 <= 1'b0;
      vvv_d_sva_10_30_0 <= 31'b0000000000000000000000000000000;
      uuu_d_sva_10_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( det_d_and_12_cse ) begin
      det_d_sva_12_30_0 <= det_d_sva_11_30_0;
      operator_1_false_return_sva_10 <= operator_1_false_return_sva_9;
      operator_1_false_return_1_sva_10 <= operator_1_false_return_1_sva_9;
      vvv_d_sva_10_30_0 <= vvv_d_sva_9_30_0;
      uuu_d_sva_10_30_0 <= uuu_d_sva_9_30_0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_1_false_return_2_sva_2 <= 1'b0;
      if_ttt_d_sva_2_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( if_and_cse ) begin
      operator_1_false_return_2_sva_2 <= operator_1_false_return_2_sva_1;
      if_ttt_d_sva_2_30_0 <= if_ttt_d_sva_1_30_0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      FP_GEQ_32_8_lor_lpi_1_dfm_2 <= 1'b0;
      ist_req_stream_rid_slc_ist_req_stream_crt_9_0_itm_2 <= 10'b0000000000;
    end
    else if ( FP_GEQ_32_8_oelse_and_cse ) begin
      FP_GEQ_32_8_lor_lpi_1_dfm_2 <= FP_GEQ_32_8_lor_lpi_1_dfm_st;
      ist_req_stream_rid_slc_ist_req_stream_crt_9_0_itm_2 <= ist_req_stream_rid_slc_ist_req_stream_crt_9_0_itm_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      land_1_lpi_1_dfm_1_st_8 <= 1'b0;
    end
    else if ( core_wen & (~((~ mux_131_cse) | and_dcpl_4 | (~ main_stage_v_21)))
        ) begin
      land_1_lpi_1_dfm_1_st_8 <= land_1_lpi_1_dfm_1_st_7;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_23 <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_47 & main_stage_v_22) | main_stage_v_23_mx0c1)
        ) begin
      main_stage_v_23 <= ~ main_stage_v_23_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_24 <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_15 & main_stage_v_23) | main_stage_v_24_mx0c1)
        ) begin
      main_stage_v_24 <= ~ main_stage_v_24_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_1_false_return_1_sva_12 <= 1'b0;
      vv_i_slc_vvv_d_30_0_itm_2 <= 31'b0000000000000000000000000000000;
      operator_1_false_return_sva_12 <= 1'b0;
      uu_i_slc_uuu_d_30_0_itm_2 <= 31'b0000000000000000000000000000000;
      operator_1_false_return_2_sva_4 <= 1'b0;
      if_tt_i_slc_if_ttt_d_30_0_itm_2 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_799_cse ) begin
      operator_1_false_return_1_sva_12 <= operator_1_false_return_1_sva_11;
      vv_i_slc_vvv_d_30_0_itm_2 <= vv_i_slc_vvv_d_30_0_itm_1;
      operator_1_false_return_sva_12 <= operator_1_false_return_sva_11;
      uu_i_slc_uuu_d_30_0_itm_2 <= uu_i_slc_uuu_d_30_0_itm_1;
      operator_1_false_return_2_sva_4 <= operator_1_false_return_2_sva_3;
      if_tt_i_slc_if_ttt_d_30_0_itm_2 <= if_tt_i_slc_if_ttt_d_30_0_itm_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      if_land_lpi_1_dfm_1_st_2 <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_25) ) begin
      if_land_lpi_1_dfm_1_st_2 <= if_land_lpi_1_dfm_1_st_1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_25 <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_56 & main_stage_v_24) | main_stage_v_25_mx0c1)
        ) begin
      main_stage_v_25 <= ~ main_stage_v_25_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_26 <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_20 & main_stage_v_25) | main_stage_v_26_mx0c1)
        ) begin
      main_stage_v_26 <= ~ main_stage_v_26_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      if_land_lpi_1_dfm_1_st_4 <= 1'b0;
    end
    else if ( core_wen & (~ or_dcpl_34) ) begin
      if_land_lpi_1_dfm_1_st_4 <= if_land_lpi_1_dfm_1_3;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      land_1_lpi_1_dfm_1_12 <= 1'b0;
      ist_req_stream_rid_slc_ist_req_stream_crt_9_0_itm_6 <= 10'b0000000000;
      if_if_if_if_and_itm_4 <= 1'b0;
    end
    else if ( if_aelse_and_10_cse ) begin
      land_1_lpi_1_dfm_1_12 <= land_1_lpi_1_dfm_1_11;
      ist_req_stream_rid_slc_ist_req_stream_crt_9_0_itm_6 <= ist_req_stream_rid_slc_ist_req_stream_crt_9_0_itm_5;
      if_if_if_if_and_itm_4 <= if_if_if_if_and_itm_3;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_20 <= 1'b0;
    end
    else if ( core_wen & (lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_20_cse
        | main_stage_v_20_mx0c1) ) begin
      main_stage_v_20 <= ~ main_stage_v_20_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ist_req_stream_crt_sva_20_265_234 <= 32'b00000000000000000000000000000000;
      det_d_sva_10 <= 32'b00000000000000000000000000000000;
      lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_24_sva_4 <= 32'b00000000000000000000000000000000;
      uuu_d_sva_8_30_0 <= 31'b0000000000000000000000000000000;
      vvv_d_sva_8_30_0 <= 31'b0000000000000000000000000000000;
      operator_1_false_return_sva_8 <= 1'b0;
      operator_1_false_return_1_sva_8 <= 1'b0;
    end
    else if ( and_801_cse ) begin
      ist_req_stream_crt_sva_20_265_234 <= ist_req_stream_crt_sva_19_265_234;
      det_d_sva_10 <= det_d_sva_9;
      lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_24_sva_4 <= lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_24_sva_3;
      uuu_d_sva_8_30_0 <= uuu_d_sva_7_30_0;
      vvv_d_sva_8_30_0 <= vvv_d_sva_7_30_0;
      operator_1_false_return_sva_8 <= operator_1_false_return_sva_7;
      operator_1_false_return_1_sva_8 <= operator_1_false_return_1_sva_7;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      land_1_lpi_1_dfm_1_st_6 <= 1'b0;
      ist_req_stream_crt_sva_20_9_0 <= 10'b0000000000;
    end
    else if ( aelse_1_and_4_cse ) begin
      land_1_lpi_1_dfm_1_st_6 <= land_1_lpi_1_dfm_1_st_5;
      ist_req_stream_crt_sva_20_9_0 <= ist_req_stream_crt_sva_19_9_0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_19 <= 1'b0;
    end
    else if ( core_wen & (lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_19_cse
        | main_stage_v_19_mx0c1) ) begin
      main_stage_v_19 <= ~ main_stage_v_19_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_18 <= 1'b0;
    end
    else if ( core_wen & (lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_18_cse
        | main_stage_v_18_mx0c1) ) begin
      main_stage_v_18 <= ~ main_stage_v_18_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_23_sva_2 <= 32'b00000000000000000000000000000000;
      ist_req_stream_crt_sva_18_265_234 <= 32'b00000000000000000000000000000000;
      det_d_sva_8 <= 32'b00000000000000000000000000000000;
      lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_24_sva_2 <= 32'b00000000000000000000000000000000;
      uuu_d_sva_6_30_0 <= 31'b0000000000000000000000000000000;
      vvv_d_sva_6_30_0 <= 31'b0000000000000000000000000000000;
      operator_1_false_return_sva_6 <= 1'b0;
      operator_1_false_return_1_sva_6 <= 1'b0;
    end
    else if ( if_and_7_cse ) begin
      lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_23_sva_2 <= lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_23_sva_1;
      ist_req_stream_crt_sva_18_265_234 <= ist_req_stream_crt_sva_17_265_234;
      det_d_sva_8 <= det_d_sva_7;
      lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_24_sva_2 <= lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_24_sva_1;
      uuu_d_sva_6_30_0 <= uuu_d_sva_5_30_0;
      vvv_d_sva_6_30_0 <= vvv_d_sva_5_30_0;
      operator_1_false_return_sva_6 <= operator_1_false_return_sva_5;
      operator_1_false_return_1_sva_6 <= operator_1_false_return_1_sva_5;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      land_1_lpi_1_dfm_1_st_4 <= 1'b0;
      ist_req_stream_crt_sva_18_9_0 <= 10'b0000000000;
    end
    else if ( aelse_1_and_5_cse ) begin
      land_1_lpi_1_dfm_1_st_4 <= land_1_lpi_1_dfm_1_st_3;
      ist_req_stream_crt_sva_18_9_0 <= ist_req_stream_crt_sva_17_9_0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_17 <= 1'b0;
    end
    else if ( core_wen & (lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_17_cse
        | main_stage_v_17_mx0c1) ) begin
      main_stage_v_17 <= ~ main_stage_v_17_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_16 <= 1'b0;
    end
    else if ( core_wen & (lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_16_cse
        | main_stage_v_16_mx0c1) ) begin
      main_stage_v_16 <= ~ main_stage_v_16_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      land_1_lpi_1_dfm_1_st_2 <= 1'b0;
      ist_req_stream_crt_sva_16_9_0 <= 10'b0000000000;
    end
    else if ( aelse_1_and_6_cse ) begin
      land_1_lpi_1_dfm_1_st_2 <= land_1_lpi_1_dfm_1_st_1;
      ist_req_stream_crt_sva_16_9_0 <= ist_req_stream_crt_sva_15_9_0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_15 <= 1'b0;
    end
    else if ( core_wen & (lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_15_cse
        | main_stage_v_15_mx0c1) ) begin
      main_stage_v_15 <= ~ main_stage_v_15_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_14 <= 1'b0;
    end
    else if ( core_wen & (lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_14_cse
        | main_stage_v_14_mx0c1) ) begin
      main_stage_v_14 <= ~ main_stage_v_14_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ist_req_stream_crt_sva_14_265_202 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      det_d_sva_4 <= 32'b00000000000000000000000000000000;
      n_z_d_sva_10 <= 32'b00000000000000000000000000000000;
      c_z_d_sva_12 <= 32'b00000000000000000000000000000000;
      n_y_d_sva_10 <= 32'b00000000000000000000000000000000;
      c_y_d_sva_12 <= 32'b00000000000000000000000000000000;
      n_x_d_sva_10 <= 32'b00000000000000000000000000000000;
      c_x_d_sva_12 <= 32'b00000000000000000000000000000000;
      uuu_d_sva_2_30_0 <= 31'b0000000000000000000000000000000;
      vvv_d_sva_2_30_0 <= 31'b0000000000000000000000000000000;
      operator_1_false_return_sva_2 <= 1'b0;
      operator_1_false_return_1_sva_2 <= 1'b0;
    end
    else if ( and_802_cse ) begin
      ist_req_stream_crt_sva_14_265_202 <= ist_req_stream_crt_sva_13_265_202;
      det_d_sva_4 <= det_d_sva_3;
      n_z_d_sva_10 <= n_z_d_sva_9;
      c_z_d_sva_12 <= c_z_d_sva_11;
      n_y_d_sva_10 <= n_y_d_sva_9;
      c_y_d_sva_12 <= c_y_d_sva_11;
      n_x_d_sva_10 <= n_x_d_sva_9;
      c_x_d_sva_12 <= c_x_d_sva_11;
      uuu_d_sva_2_30_0 <= uuu_d_sva_1_30_0;
      vvv_d_sva_2_30_0 <= vvv_d_sva_1_30_0;
      operator_1_false_return_sva_2 <= ccs_lp_piped_fp_add_23_8_0_cmp_3_a_core_31;
      operator_1_false_return_1_sva_2 <= ccs_lp_piped_fp_add_23_8_0_cmp_3_b_core_31;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      fp_arelb_32_8_return_0_sva <= 1'b0;
      FP_LEQ_32_8_arelb_1_sva <= 1'b0;
    end
    else if ( FP_LEQ_32_8_arelb_and_cse ) begin
      fp_arelb_32_8_return_0_sva <= ccs_fp_cmp_23_8_0_out_6;
      FP_LEQ_32_8_arelb_1_sva <= ccs_fp_cmp_23_8_0_out_7;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      land_lpi_1_dfm_2 <= 1'b0;
      ist_req_stream_crt_sva_14_9_0 <= 10'b0000000000;
    end
    else if ( aelse_and_cse ) begin
      land_lpi_1_dfm_2 <= land_lpi_1_dfm_1;
      ist_req_stream_crt_sva_14_9_0 <= ist_req_stream_crt_sva_13_9_0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_13 <= 1'b0;
    end
    else if ( core_wen & (lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_13_cse
        | main_stage_v_13_mx0c1) ) begin
      main_stage_v_13 <= ~ main_stage_v_13_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_12 <= 1'b0;
    end
    else if ( core_wen & (lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_12_cse
        | main_stage_v_12_mx0c1) ) begin
      main_stage_v_12 <= ~ main_stage_v_12_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      det_d_sva_2 <= 32'b00000000000000000000000000000000;
      ist_req_stream_crt_sva_12_265_202 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      n_x_d_sva_8 <= 32'b00000000000000000000000000000000;
      n_y_d_sva_8 <= 32'b00000000000000000000000000000000;
      n_z_d_sva_8 <= 32'b00000000000000000000000000000000;
      c_x_d_sva_10 <= 32'b00000000000000000000000000000000;
      c_y_d_sva_10 <= 32'b00000000000000000000000000000000;
      c_z_d_sva_10 <= 32'b00000000000000000000000000000000;
      ist_req_stream_crt_sva_12_9_0 <= 10'b0000000000;
    end
    else if ( det_d_and_3_cse ) begin
      det_d_sva_2 <= det_d_sva_1;
      ist_req_stream_crt_sva_12_265_202 <= ist_req_stream_crt_sva_11_265_202;
      n_x_d_sva_8 <= n_x_d_sva_7;
      n_y_d_sva_8 <= n_y_d_sva_7;
      n_z_d_sva_8 <= n_z_d_sva_7;
      c_x_d_sva_10 <= c_x_d_sva_9;
      c_y_d_sva_10 <= c_y_d_sva_9;
      c_z_d_sva_10 <= c_z_d_sva_9;
      ist_req_stream_crt_sva_12_9_0 <= ist_req_stream_crt_sva_11_9_0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_11 <= 1'b0;
    end
    else if ( core_wen & (lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_11_cse
        | main_stage_v_11_mx0c1) ) begin
      main_stage_v_11 <= ~ main_stage_v_11_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_10 <= 1'b0;
    end
    else if ( core_wen & (lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_10_cse
        | main_stage_v_10_mx0c1) ) begin
      main_stage_v_10 <= ~ main_stage_v_10_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_20_sva_2 <= 32'b00000000000000000000000000000000;
      lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_17_sva_2 <= 32'b00000000000000000000000000000000;
      ist_req_stream_crt_sva_10_265_202 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      n_x_d_sva_6 <= 32'b00000000000000000000000000000000;
      n_y_d_sva_6 <= 32'b00000000000000000000000000000000;
      n_z_d_sva_6 <= 32'b00000000000000000000000000000000;
      c_x_d_sva_8 <= 32'b00000000000000000000000000000000;
      c_y_d_sva_8 <= 32'b00000000000000000000000000000000;
      c_z_d_sva_8 <= 32'b00000000000000000000000000000000;
      ist_req_stream_crt_sva_10_9_0 <= 10'b0000000000;
    end
    else if ( and_660_cse ) begin
      lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_20_sva_2 <= lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_20_sva_1;
      lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_17_sva_2 <= lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_17_sva_1;
      ist_req_stream_crt_sva_10_265_202 <= ist_req_stream_crt_sva_9_265_202;
      n_x_d_sva_6 <= n_x_d_sva_5;
      n_y_d_sva_6 <= n_y_d_sva_5;
      n_z_d_sva_6 <= n_z_d_sva_5;
      c_x_d_sva_8 <= c_x_d_sva_7;
      c_y_d_sva_8 <= c_y_d_sva_7;
      c_z_d_sva_8 <= c_z_d_sva_7;
      ist_req_stream_crt_sva_10_9_0 <= ist_req_stream_crt_sva_9_9_0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_9 <= 1'b0;
    end
    else if ( core_wen & (lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_9_cse
        | main_stage_v_9_mx0c1) ) begin
      main_stage_v_9 <= ~ main_stage_v_9_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_8 <= 1'b0;
    end
    else if ( core_wen & (lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_8_cse
        | main_stage_v_8_mx0c1) ) begin
      main_stage_v_8 <= ~ main_stage_v_8_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_14_sva_2 <= 32'b00000000000000000000000000000000;
      ist_req_stream_crt_sva_8_265_202 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      n_x_d_sva_4 <= 32'b00000000000000000000000000000000;
      n_y_d_sva_4 <= 32'b00000000000000000000000000000000;
      n_z_d_sva_4 <= 32'b00000000000000000000000000000000;
      c_x_d_sva_6 <= 32'b00000000000000000000000000000000;
      c_y_d_sva_6 <= 32'b00000000000000000000000000000000;
      c_z_d_sva_6 <= 32'b00000000000000000000000000000000;
      ist_req_stream_crt_sva_8_9_0 <= 10'b0000000000;
    end
    else if ( and_664_cse ) begin
      lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_14_sva_2 <= lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_14_sva_1;
      ist_req_stream_crt_sva_8_265_202 <= ist_req_stream_crt_sva_7_265_202;
      n_x_d_sva_4 <= n_x_d_sva_3;
      n_y_d_sva_4 <= n_y_d_sva_3;
      n_z_d_sva_4 <= n_z_d_sva_3;
      c_x_d_sva_6 <= c_x_d_sva_5;
      c_y_d_sva_6 <= c_y_d_sva_5;
      c_z_d_sva_6 <= c_z_d_sva_5;
      ist_req_stream_crt_sva_8_9_0 <= ist_req_stream_crt_sva_7_9_0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_7 <= 1'b0;
    end
    else if ( core_wen & (lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_7_cse
        | main_stage_v_7_mx0c1) ) begin
      main_stage_v_7 <= ~ main_stage_v_7_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_6 <= 1'b0;
    end
    else if ( core_wen & (lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_6_cse
        | main_stage_v_6_mx0c1) ) begin
      main_stage_v_6 <= ~ main_stage_v_6_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ist_req_stream_crt_sva_6_553_362 <= 192'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      ist_req_stream_crt_sva_6_265_202 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      n_x_d_sva_2 <= 32'b00000000000000000000000000000000;
      n_y_d_sva_2 <= 32'b00000000000000000000000000000000;
      n_z_d_sva_2 <= 32'b00000000000000000000000000000000;
      c_x_d_sva_4 <= 32'b00000000000000000000000000000000;
      c_y_d_sva_4 <= 32'b00000000000000000000000000000000;
      c_z_d_sva_4 <= 32'b00000000000000000000000000000000;
      ist_req_stream_crt_sva_6_9_0 <= 10'b0000000000;
    end
    else if ( and_667_cse ) begin
      ist_req_stream_crt_sva_6_553_362 <= ist_req_stream_crt_sva_5_553_362;
      ist_req_stream_crt_sva_6_265_202 <= ist_req_stream_crt_sva_5_265_202;
      n_x_d_sva_2 <= n_x_d_sva_1;
      n_y_d_sva_2 <= n_y_d_sva_1;
      n_z_d_sva_2 <= n_z_d_sva_1;
      c_x_d_sva_4 <= c_x_d_sva_3;
      c_y_d_sva_4 <= c_y_d_sva_3;
      c_z_d_sva_4 <= c_z_d_sva_3;
      ist_req_stream_crt_sva_6_9_0 <= ist_req_stream_crt_sva_5_9_0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_5 <= 1'b0;
    end
    else if ( core_wen & (lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_5_cse
        | main_stage_v_5_mx0c1) ) begin
      main_stage_v_5 <= ~ main_stage_v_5_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_4 <= 1'b0;
    end
    else if ( core_wen & (lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_4_cse
        | main_stage_v_4_mx0c1) ) begin
      main_stage_v_4 <= ~ main_stage_v_4_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ist_req_stream_crt_sva_4_265_106 <= 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      ist_req_stream_crt_sva_4_553_362 <= 192'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      c_x_d_sva_2 <= 32'b00000000000000000000000000000000;
      c_y_d_sva_2 <= 32'b00000000000000000000000000000000;
      c_z_d_sva_2 <= 32'b00000000000000000000000000000000;
      ist_req_stream_crt_sva_4_9_0 <= 10'b0000000000;
    end
    else if ( and_670_cse ) begin
      ist_req_stream_crt_sva_4_265_106 <= ist_req_stream_crt_sva_3_265_106;
      ist_req_stream_crt_sva_4_553_362 <= ist_req_stream_crt_sva_3_553_362;
      c_x_d_sva_2 <= c_x_d_sva_1;
      c_y_d_sva_2 <= c_y_d_sva_1;
      c_z_d_sva_2 <= c_z_d_sva_1;
      ist_req_stream_crt_sva_4_9_0 <= ist_req_stream_crt_sva_3_9_0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_3 <= 1'b0;
    end
    else if ( core_wen & (lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_3_cse
        | main_stage_v_3_mx0c1) ) begin
      main_stage_v_3 <= ~ main_stage_v_3_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_2 <= 1'b0;
    end
    else if ( core_wen & (lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_2_cse
        | main_stage_v_2_mx0c1) ) begin
      main_stage_v_2 <= ~ main_stage_v_2_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ist_req_stream_crt_sva_2_265_106 <= 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      ist_req_stream_crt_sva_2_553_362 <= 192'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      ist_req_stream_crt_sva_2_9_0 <= 10'b0000000000;
    end
    else if ( and_673_cse ) begin
      ist_req_stream_crt_sva_2_265_106 <= ist_req_stream_crt_sva_1_265_106;
      ist_req_stream_crt_sva_2_553_362 <= ist_req_stream_crt_sva_1_553_362;
      ist_req_stream_crt_sva_2_9_0 <= ist_req_stream_crt_sva_1_9_0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      main_stage_v_1 <= 1'b0;
    end
    else if ( core_wen & (lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_lp_piped_fp_mult_AC_RND_CONV_0_32_8_rnd_and_1_cse
        | main_stage_v_1_mx0c1) ) begin
      main_stage_v_1 <= ~ main_stage_v_1_mx0c1;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      det_d_sva_11_30_0 <= 31'b0000000000000000000000000000000;
      uuu_d_sva_9_30_0 <= 31'b0000000000000000000000000000000;
      vvv_d_sva_9_30_0 <= 31'b0000000000000000000000000000000;
      operator_1_false_return_sva_9 <= 1'b0;
      operator_1_false_return_1_sva_9 <= 1'b0;
    end
    else if ( det_d_and_15_cse ) begin
      det_d_sva_11_30_0 <= det_d_sva_10[30:0];
      uuu_d_sva_9_30_0 <= uuu_d_sva_8_30_0;
      vvv_d_sva_9_30_0 <= vvv_d_sva_8_30_0;
      operator_1_false_return_sva_9 <= operator_1_false_return_sva_8;
      operator_1_false_return_1_sva_9 <= operator_1_false_return_1_sva_8;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      if_ttt_d_sva_1_30_0 <= 31'b0000000000000000000000000000000;
      operator_1_false_return_2_sva_1 <= 1'b0;
    end
    else if ( if_ttt_d_and_2_cse ) begin
      if_ttt_d_sva_1_30_0 <= ccs_lp_piped_fp_add_23_8_0_cmp_1_z_mxwt[30:0];
      operator_1_false_return_2_sva_1 <= operator_1_false_return_2_sva_mx0w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      land_1_lpi_1_dfm_1_st_7 <= 1'b0;
      ist_req_stream_rid_slc_ist_req_stream_crt_9_0_itm_1 <= 10'b0000000000;
    end
    else if ( det_d_and_4_cse ) begin
      land_1_lpi_1_dfm_1_st_7 <= land_1_lpi_1_dfm_1_st_6;
      ist_req_stream_rid_slc_ist_req_stream_crt_9_0_itm_1 <= ist_req_stream_crt_sva_20_9_0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      operator_1_false_return_sva_11 <= 1'b0;
      operator_1_false_return_1_sva_11 <= 1'b0;
      operator_1_false_return_2_sva_3 <= 1'b0;
      if_tt_i_slc_if_ttt_d_30_0_itm_1 <= 31'b0000000000000000000000000000000;
      uu_i_slc_uuu_d_30_0_itm_1 <= 31'b0000000000000000000000000000000;
      vv_i_slc_vvv_d_30_0_itm_1 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_803_cse ) begin
      operator_1_false_return_sva_11 <= operator_1_false_return_sva_10;
      operator_1_false_return_1_sva_11 <= operator_1_false_return_1_sva_10;
      operator_1_false_return_2_sva_3 <= operator_1_false_return_2_sva_2;
      if_tt_i_slc_if_ttt_d_30_0_itm_1 <= if_ttt_d_sva_2_30_0;
      uu_i_slc_uuu_d_30_0_itm_1 <= uuu_d_sva_10_30_0;
      vv_i_slc_vvv_d_30_0_itm_1 <= vvv_d_sva_10_30_0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      land_1_lpi_1_dfm_1_st_9 <= 1'b0;
      if_if_if_if_and_itm_1 <= 1'b0;
      ist_req_stream_rid_slc_ist_req_stream_crt_9_0_itm_3 <= 10'b0000000000;
    end
    else if ( aelse_1_and_25_cse ) begin
      land_1_lpi_1_dfm_1_st_9 <= land_1_lpi_1_dfm_1_st_8;
      if_if_if_if_and_itm_1 <= if_land_lpi_1_dfm_2 & FP_GEQ_32_8_lor_lpi_1_dfm_2
          & land_1_lpi_1_dfm_1_st_8;
      ist_req_stream_rid_slc_ist_req_stream_crt_9_0_itm_3 <= ist_req_stream_rid_slc_ist_req_stream_crt_9_0_itm_2;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      if_land_lpi_1_dfm_1_st_1 <= 1'b0;
    end
    else if ( core_wen & ((and_dcpl_15 & land_1_lpi_1_dfm_1_st_8) | and_dcpl_110)
        & mux_tmp_66 ) begin
      if_land_lpi_1_dfm_1_st_1 <= MUX_s_1_2_2(if_land_lpi_1_dfm_1_mx0w0, if_land_lpi_1_dfm_1_st,
          and_dcpl_110);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      land_1_lpi_1_dfm_1_11 <= 1'b0;
      if_land_lpi_1_dfm_1_3 <= 1'b0;
      if_if_if_if_and_itm_3 <= 1'b0;
      ist_req_stream_rid_slc_ist_req_stream_crt_9_0_itm_5 <= 10'b0000000000;
    end
    else if ( aelse_1_and_26_cse ) begin
      land_1_lpi_1_dfm_1_11 <= land_1_lpi_1_dfm_1_10;
      if_land_lpi_1_dfm_1_3 <= if_land_lpi_1_dfm_1_st_2;
      if_if_if_if_and_itm_3 <= if_if_if_if_and_itm_2;
      ist_req_stream_rid_slc_ist_req_stream_crt_9_0_itm_5 <= ist_req_stream_rid_slc_ist_req_stream_crt_9_0_itm_4;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ist_req_stream_crt_sva_13_265_202 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      n_x_d_sva_9 <= 32'b00000000000000000000000000000000;
      n_y_d_sva_9 <= 32'b00000000000000000000000000000000;
      n_z_d_sva_9 <= 32'b00000000000000000000000000000000;
      c_x_d_sva_11 <= 32'b00000000000000000000000000000000;
      c_y_d_sva_11 <= 32'b00000000000000000000000000000000;
      c_z_d_sva_11 <= 32'b00000000000000000000000000000000;
      det_d_sva_3 <= 32'b00000000000000000000000000000000;
      uuu_d_sva_1_30_0 <= 31'b0000000000000000000000000000000;
      vvv_d_sva_1_30_0 <= 31'b0000000000000000000000000000000;
    end
    else if ( and_805_cse ) begin
      ist_req_stream_crt_sva_13_265_202 <= ist_req_stream_crt_sva_12_265_202;
      n_x_d_sva_9 <= n_x_d_sva_8;
      n_y_d_sva_9 <= n_y_d_sva_8;
      n_z_d_sva_9 <= n_z_d_sva_8;
      c_x_d_sva_11 <= c_x_d_sva_10;
      c_y_d_sva_11 <= c_y_d_sva_10;
      c_z_d_sva_11 <= c_z_d_sva_10;
      det_d_sva_3 <= det_d_sva_2;
      uuu_d_sva_1_30_0 <= ccs_lp_piped_fp_add_23_8_0_cmp_6_z_mxwt[30:0];
      vvv_d_sva_1_30_0 <= ccs_lp_piped_fp_add_23_8_0_cmp_4_z_mxwt[30:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ist_req_stream_crt_sva_19_265_234 <= 32'b00000000000000000000000000000000;
      det_d_sva_9 <= 32'b00000000000000000000000000000000;
      lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_24_sva_3 <= 32'b00000000000000000000000000000000;
      uuu_d_sva_7_30_0 <= 31'b0000000000000000000000000000000;
      vvv_d_sva_7_30_0 <= 31'b0000000000000000000000000000000;
      operator_1_false_return_sva_7 <= 1'b0;
      operator_1_false_return_1_sva_7 <= 1'b0;
    end
    else if ( and_806_cse ) begin
      ist_req_stream_crt_sva_19_265_234 <= ist_req_stream_crt_sva_18_265_234;
      det_d_sva_9 <= det_d_sva_8;
      lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_24_sva_3 <= lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_24_sva_2;
      uuu_d_sva_7_30_0 <= uuu_d_sva_6_30_0;
      vvv_d_sva_7_30_0 <= vvv_d_sva_6_30_0;
      operator_1_false_return_sva_7 <= operator_1_false_return_sva_6;
      operator_1_false_return_1_sva_7 <= operator_1_false_return_1_sva_6;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ist_req_stream_crt_sva_5_553_362 <= 192'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      ist_req_stream_crt_sva_5_265_202 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      n_x_d_sva_1 <= 32'b00000000000000000000000000000000;
      n_y_d_sva_1 <= 32'b00000000000000000000000000000000;
      n_z_d_sva_1 <= 32'b00000000000000000000000000000000;
      c_x_d_sva_3 <= 32'b00000000000000000000000000000000;
      c_y_d_sva_3 <= 32'b00000000000000000000000000000000;
      c_z_d_sva_3 <= 32'b00000000000000000000000000000000;
      ist_req_stream_crt_sva_5_9_0 <= 10'b0000000000;
    end
    else if ( and_679_cse ) begin
      ist_req_stream_crt_sva_5_553_362 <= ist_req_stream_crt_sva_4_553_362;
      ist_req_stream_crt_sva_5_265_202 <= ist_req_stream_crt_sva_4_265_106[159:96];
      n_x_d_sva_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_z_mxwt;
      n_y_d_sva_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_17_z_mxwt;
      n_z_d_sva_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_16_z_mxwt;
      c_x_d_sva_3 <= c_x_d_sva_2;
      c_y_d_sva_3 <= c_y_d_sva_2;
      c_z_d_sva_3 <= c_z_d_sva_2;
      ist_req_stream_crt_sva_5_9_0 <= ist_req_stream_crt_sva_4_9_0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ist_req_stream_crt_sva_3_265_106 <= 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      ist_req_stream_crt_sva_3_553_362 <= 192'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      c_x_d_sva_1 <= 32'b00000000000000000000000000000000;
      c_y_d_sva_1 <= 32'b00000000000000000000000000000000;
      c_z_d_sva_1 <= 32'b00000000000000000000000000000000;
      ist_req_stream_crt_sva_3_9_0 <= 10'b0000000000;
    end
    else if ( and_680_cse ) begin
      ist_req_stream_crt_sva_3_265_106 <= ist_req_stream_crt_sva_2_265_106;
      ist_req_stream_crt_sva_3_553_362 <= ist_req_stream_crt_sva_2_553_362;
      c_x_d_sva_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_15_z_mxwt;
      c_y_d_sva_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_14_z_mxwt;
      c_z_d_sva_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_13_z_mxwt;
      ist_req_stream_crt_sva_3_9_0 <= ist_req_stream_crt_sva_2_9_0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ist_req_stream_crt_sva_1_265_106 <= 160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      ist_req_stream_crt_sva_1_553_362 <= 192'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      ist_req_stream_crt_sva_1_9_0 <= 10'b0000000000;
    end
    else if ( and_681_cse ) begin
      ist_req_stream_crt_sva_1_265_106 <= ist_req_stream_rsci_idat_mxwt[265:106];
      ist_req_stream_crt_sva_1_553_362 <= ist_req_stream_rsci_idat_mxwt[553:362];
      ist_req_stream_crt_sva_1_9_0 <= ist_req_stream_rsci_idat_mxwt[9:0];
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_14_sva_1 <= 32'b00000000000000000000000000000000;
      ist_req_stream_crt_sva_7_265_202 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      n_x_d_sva_3 <= 32'b00000000000000000000000000000000;
      n_y_d_sva_3 <= 32'b00000000000000000000000000000000;
      n_z_d_sva_3 <= 32'b00000000000000000000000000000000;
      c_x_d_sva_5 <= 32'b00000000000000000000000000000000;
      c_y_d_sva_5 <= 32'b00000000000000000000000000000000;
      c_z_d_sva_5 <= 32'b00000000000000000000000000000000;
      ist_req_stream_crt_sva_7_9_0 <= 10'b0000000000;
    end
    else if ( and_682_cse ) begin
      lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_14_sva_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_15_z_mxwt;
      ist_req_stream_crt_sva_7_265_202 <= ist_req_stream_crt_sva_6_265_202;
      n_x_d_sva_3 <= n_x_d_sva_2;
      n_y_d_sva_3 <= n_y_d_sva_2;
      n_z_d_sva_3 <= n_z_d_sva_2;
      c_x_d_sva_5 <= c_x_d_sva_4;
      c_y_d_sva_5 <= c_y_d_sva_4;
      c_z_d_sva_5 <= c_z_d_sva_4;
      ist_req_stream_crt_sva_7_9_0 <= ist_req_stream_crt_sva_6_9_0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      det_d_sva_1 <= 32'b00000000000000000000000000000000;
      ist_req_stream_crt_sva_11_265_202 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      n_x_d_sva_7 <= 32'b00000000000000000000000000000000;
      n_y_d_sva_7 <= 32'b00000000000000000000000000000000;
      n_z_d_sva_7 <= 32'b00000000000000000000000000000000;
      c_x_d_sva_9 <= 32'b00000000000000000000000000000000;
      c_y_d_sva_9 <= 32'b00000000000000000000000000000000;
      c_z_d_sva_9 <= 32'b00000000000000000000000000000000;
      ist_req_stream_crt_sva_11_9_0 <= 10'b0000000000;
    end
    else if ( det_d_and_7_cse ) begin
      det_d_sva_1 <= ccs_lp_piped_fp_add_23_8_0_cmp_8_z_mxwt;
      ist_req_stream_crt_sva_11_265_202 <= ist_req_stream_crt_sva_10_265_202;
      n_x_d_sva_7 <= n_x_d_sva_6;
      n_y_d_sva_7 <= n_y_d_sva_6;
      n_z_d_sva_7 <= n_z_d_sva_6;
      c_x_d_sva_9 <= c_x_d_sva_8;
      c_y_d_sva_9 <= c_y_d_sva_8;
      c_z_d_sva_9 <= c_z_d_sva_8;
      ist_req_stream_crt_sva_11_9_0 <= ist_req_stream_crt_sva_10_9_0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_17_sva_1 <= 32'b00000000000000000000000000000000;
      lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_20_sva_1 <= 32'b00000000000000000000000000000000;
      ist_req_stream_crt_sva_9_265_202 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      n_x_d_sva_5 <= 32'b00000000000000000000000000000000;
      n_y_d_sva_5 <= 32'b00000000000000000000000000000000;
      n_z_d_sva_5 <= 32'b00000000000000000000000000000000;
      c_x_d_sva_7 <= 32'b00000000000000000000000000000000;
      c_y_d_sva_7 <= 32'b00000000000000000000000000000000;
      c_z_d_sva_7 <= 32'b00000000000000000000000000000000;
      ist_req_stream_crt_sva_9_9_0 <= 10'b0000000000;
    end
    else if ( and_683_cse ) begin
      lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_17_sva_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_12_z_mxwt;
      lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_20_sva_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_9_z_mxwt;
      ist_req_stream_crt_sva_9_265_202 <= ist_req_stream_crt_sva_8_265_202;
      n_x_d_sva_5 <= n_x_d_sva_4;
      n_y_d_sva_5 <= n_y_d_sva_4;
      n_z_d_sva_5 <= n_z_d_sva_4;
      c_x_d_sva_7 <= c_x_d_sva_6;
      c_y_d_sva_7 <= c_y_d_sva_6;
      c_z_d_sva_7 <= c_z_d_sva_6;
      ist_req_stream_crt_sva_9_9_0 <= ist_req_stream_crt_sva_8_9_0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      land_lpi_1_dfm_1 <= 1'b0;
      ist_req_stream_crt_sva_13_9_0 <= 10'b0000000000;
    end
    else if ( aelse_and_2_cse ) begin
      land_lpi_1_dfm_1 <= nor_105_cse;
      ist_req_stream_crt_sva_13_9_0 <= ist_req_stream_crt_sva_12_9_0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_23_sva_1 <= 32'b00000000000000000000000000000000;
      ist_req_stream_crt_sva_17_265_234 <= 32'b00000000000000000000000000000000;
      det_d_sva_7 <= 32'b00000000000000000000000000000000;
      lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_24_sva_1 <= 32'b00000000000000000000000000000000;
      uuu_d_sva_5_30_0 <= 31'b0000000000000000000000000000000;
      vvv_d_sva_5_30_0 <= 31'b0000000000000000000000000000000;
      operator_1_false_return_sva_5 <= 1'b0;
      operator_1_false_return_1_sva_5 <= 1'b0;
    end
    else if ( if_and_10_cse ) begin
      lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_23_sva_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_6_z_mxwt;
      ist_req_stream_crt_sva_17_265_234 <= ist_req_stream_crt_sva_16_265_234;
      det_d_sva_7 <= det_d_sva_6;
      lp_piped_fp_mult_AC_RND_CONV_0_32_8_return_d_24_sva_1 <= ccs_lp_piped_fp_mult_23_8_0_cmp_5_z_mxwt;
      uuu_d_sva_5_30_0 <= uuu_d_sva_4_30_0;
      vvv_d_sva_5_30_0 <= vvv_d_sva_4_30_0;
      operator_1_false_return_sva_5 <= operator_1_false_return_sva_4;
      operator_1_false_return_1_sva_5 <= operator_1_false_return_1_sva_4;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      land_1_lpi_1_dfm_1_st_5 <= 1'b0;
      ist_req_stream_crt_sva_19_9_0 <= 10'b0000000000;
    end
    else if ( aelse_1_and_11_cse ) begin
      land_1_lpi_1_dfm_1_st_5 <= land_1_lpi_1_dfm_1_st_4;
      ist_req_stream_crt_sva_19_9_0 <= ist_req_stream_crt_sva_18_9_0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      land_1_lpi_1_dfm_1_st_3 <= 1'b0;
      ist_req_stream_crt_sva_17_9_0 <= 10'b0000000000;
    end
    else if ( aelse_1_and_12_cse ) begin
      land_1_lpi_1_dfm_1_st_3 <= land_1_lpi_1_dfm_1_st_2;
      ist_req_stream_crt_sva_17_9_0 <= ist_req_stream_crt_sva_16_9_0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      land_1_lpi_1_dfm_1_st_1 <= 1'b0;
      ist_req_stream_crt_sva_15_9_0 <= 10'b0000000000;
    end
    else if ( aelse_1_and_13_cse ) begin
      land_1_lpi_1_dfm_1_st_1 <= FP_LEQ_32_8_FP_LEQ_32_8_or_cse & land_lpi_1_dfm_2;
      ist_req_stream_crt_sva_15_9_0 <= ist_req_stream_crt_sva_14_9_0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      if_land_lpi_1_dfm_1_st <= 1'b0;
    end
    else if ( core_wen & (~((~(land_1_lpi_1_dfm_1_st_8 & main_stage_v_22)) | (fsm_output[0])))
        & (~ mux_104_nl) ) begin
      if_land_lpi_1_dfm_1_st <= if_land_lpi_1_dfm_1_mx0w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      land_1_lpi_1_dfm_1_10 <= 1'b0;
      if_if_if_if_and_itm_2 <= 1'b0;
      ist_req_stream_rid_slc_ist_req_stream_crt_9_0_itm_4 <= 10'b0000000000;
    end
    else if ( aelse_1_and_28_cse ) begin
      land_1_lpi_1_dfm_1_10 <= land_1_lpi_1_dfm_1_st_9;
      if_if_if_if_and_itm_2 <= if_if_if_if_and_itm_1;
      ist_req_stream_rid_slc_ist_req_stream_crt_9_0_itm_4 <= ist_req_stream_rid_slc_ist_req_stream_crt_9_0_itm_3;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      FP_GEQ_32_8_lor_lpi_1_dfm_st <= 1'b0;
    end
    else if ( core_wen & land_1_lpi_1_dfm_1_st_6 & and_15_tmp ) begin
      FP_GEQ_32_8_lor_lpi_1_dfm_st <= or_620_cse;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ist_req_stream_crt_sva_16_265_234 <= 32'b00000000000000000000000000000000;
      det_d_sva_6 <= 32'b00000000000000000000000000000000;
      uuu_d_sva_4_30_0 <= 31'b0000000000000000000000000000000;
      vvv_d_sva_4_30_0 <= 31'b0000000000000000000000000000000;
      operator_1_false_return_sva_4 <= 1'b0;
      operator_1_false_return_1_sva_4 <= 1'b0;
    end
    else if ( and_815_cse ) begin
      ist_req_stream_crt_sva_16_265_234 <= ist_req_stream_crt_sva_15_265_234;
      det_d_sva_6 <= det_d_sva_5;
      uuu_d_sva_4_30_0 <= uuu_d_sva_3_30_0;
      vvv_d_sva_4_30_0 <= vvv_d_sva_3_30_0;
      operator_1_false_return_sva_4 <= operator_1_false_return_sva_3;
      operator_1_false_return_1_sva_4 <= operator_1_false_return_1_sva_3;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      ist_req_stream_crt_sva_15_265_234 <= 32'b00000000000000000000000000000000;
      det_d_sva_5 <= 32'b00000000000000000000000000000000;
      uuu_d_sva_3_30_0 <= 31'b0000000000000000000000000000000;
      vvv_d_sva_3_30_0 <= 31'b0000000000000000000000000000000;
      operator_1_false_return_sva_3 <= 1'b0;
      operator_1_false_return_1_sva_3 <= 1'b0;
    end
    else if ( and_816_cse ) begin
      ist_req_stream_crt_sva_15_265_234 <= ist_req_stream_crt_sva_14_265_202[63:32];
      det_d_sva_5 <= det_d_sva_4;
      uuu_d_sva_3_30_0 <= uuu_d_sva_2_30_0;
      vvv_d_sva_3_30_0 <= vvv_d_sva_2_30_0;
      operator_1_false_return_sva_3 <= operator_1_false_return_sva_2;
      operator_1_false_return_1_sva_3 <= operator_1_false_return_1_sva_2;
    end
  end
  assign or_575_nl = (~ main_stage_v_21) | land_1_lpi_1_dfm_1_st_7;
  assign mux_99_nl = MUX_s_1_2_2((~ nand_tmp_3), or_tmp_15, or_575_nl);
  assign mux_98_nl = MUX_s_1_2_2(mux_tmp_21, mux_tmp_20, and_761_cse);
  assign mux_100_nl = MUX_s_1_2_2(mux_99_nl, mux_98_nl, main_stage_v_26);
  assign and_762_nl = main_stage_v_25 & if_land_lpi_1_dfm_1_3 & land_1_lpi_1_dfm_1_11;
  assign mux_101_nl = MUX_s_1_2_2(mux_100_nl, mux_tmp_22, and_762_nl);
  assign mux_102_nl = MUX_s_1_2_2(mux_101_nl, mux_tmp_22, and_763_cse);
  assign mux_103_nl = MUX_s_1_2_2(mux_tmp_22, mux_102_nl, and_764_cse);
  assign mux_104_nl = MUX_s_1_2_2(and_743_cse, mux_103_nl, nand_217_cse);

  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    init
// ------------------------------------------------------------------


module init (
  clk, arst_n, init_req_stream_rsc_dat, init_req_stream_rsc_vld, init_req_stream_rsc_rdy,
      trv_req_stream_rsc_dat, trv_req_stream_rsc_vld, trv_req_stream_rsc_rdy
);
  input clk;
  input arst_n;
  input [361:0] init_req_stream_rsc_dat;
  input init_req_stream_rsc_vld;
  output init_req_stream_rsc_rdy;
  output [457:0] trv_req_stream_rsc_dat;
  output trv_req_stream_rsc_vld;
  input trv_req_stream_rsc_rdy;



  // Interconnect Declarations for Component Instantiations 
  init_core init_core_inst (
      .clk(clk),
      .arst_n(arst_n),
      .init_req_stream_rsc_dat(init_req_stream_rsc_dat),
      .init_req_stream_rsc_vld(init_req_stream_rsc_vld),
      .init_req_stream_rsc_rdy(init_req_stream_rsc_rdy),
      .trv_req_stream_rsc_dat(trv_req_stream_rsc_dat),
      .trv_req_stream_rsc_vld(trv_req_stream_rsc_vld),
      .trv_req_stream_rsc_rdy(trv_req_stream_rsc_rdy)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    bbox
// ------------------------------------------------------------------


module bbox (
  clk, arst_n, bbox_req_stream_rsc_dat, bbox_req_stream_rsc_vld, bbox_req_stream_rsc_rdy,
      bbox_resp_stream_rsc_dat, bbox_resp_stream_rsc_vld, bbox_resp_stream_rsc_rdy
);
  input clk;
  input arst_n;
  input [385:0] bbox_req_stream_rsc_dat;
  input bbox_req_stream_rsc_vld;
  output bbox_req_stream_rsc_rdy;
  output [204:0] bbox_resp_stream_rsc_dat;
  output bbox_resp_stream_rsc_vld;
  input bbox_resp_stream_rsc_rdy;



  // Interconnect Declarations for Component Instantiations 
  bbox_core bbox_core_inst (
      .clk(clk),
      .arst_n(arst_n),
      .bbox_req_stream_rsc_dat(bbox_req_stream_rsc_dat),
      .bbox_req_stream_rsc_vld(bbox_req_stream_rsc_vld),
      .bbox_req_stream_rsc_rdy(bbox_req_stream_rsc_rdy),
      .bbox_resp_stream_rsc_dat(bbox_resp_stream_rsc_dat),
      .bbox_resp_stream_rsc_vld(bbox_resp_stream_rsc_vld),
      .bbox_resp_stream_rsc_rdy(bbox_resp_stream_rsc_rdy)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    ist
// ------------------------------------------------------------------


module ist (
  clk, arst_n, ist_req_stream_rsc_dat, ist_req_stream_rsc_vld, ist_req_stream_rsc_rdy,
      ist_resp_stream_rsc_dat, ist_resp_stream_rsc_vld, ist_resp_stream_rsc_rdy
);
  input clk;
  input arst_n;
  input [553:0] ist_req_stream_rsc_dat;
  input ist_req_stream_rsc_vld;
  output ist_req_stream_rsc_rdy;
  output [106:0] ist_resp_stream_rsc_dat;
  output ist_resp_stream_rsc_vld;
  input ist_resp_stream_rsc_rdy;



  // Interconnect Declarations for Component Instantiations 
  ist_core ist_core_inst (
      .clk(clk),
      .arst_n(arst_n),
      .ist_req_stream_rsc_dat(ist_req_stream_rsc_dat),
      .ist_req_stream_rsc_vld(ist_req_stream_rsc_vld),
      .ist_req_stream_rsc_rdy(ist_req_stream_rsc_rdy),
      .ist_resp_stream_rsc_dat(ist_resp_stream_rsc_dat),
      .ist_resp_stream_rsc_vld(ist_resp_stream_rsc_vld),
      .ist_resp_stream_rsc_rdy(ist_resp_stream_rsc_rdy)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    rtcore_struct
// ------------------------------------------------------------------


module rtcore_struct (
  clk, arst_n, init_req_stream_rsc_dat_d, init_req_stream_rsc_dat_d_1, init_req_stream_rsc_dat_d_2,
      init_req_stream_rsc_dat_d_3, init_req_stream_rsc_dat_d_4, init_req_stream_rsc_dat_d_5,
      init_req_stream_rsc_dat_d_6, init_req_stream_rsc_dat_d_7, init_req_stream_rsc_dat_d_8,
      init_req_stream_rsc_dat_d_9, init_req_stream_rsc_dat_d_10, init_req_stream_rsc_dat_rid,
      init_req_stream_rsc_vld, init_req_stream_rsc_rdy, bbox_req_stream_rsc_dat_z_max,
      bbox_req_stream_rsc_dat_z_min, bbox_req_stream_rsc_dat_y_max, bbox_req_stream_rsc_dat_y_min,
      bbox_req_stream_rsc_dat_x_max, bbox_req_stream_rsc_dat_x_min, bbox_req_stream_rsc_dat_z_max_1,
      bbox_req_stream_rsc_dat_z_min_1, bbox_req_stream_rsc_dat_y_max_1, bbox_req_stream_rsc_dat_y_min_1,
      bbox_req_stream_rsc_dat_x_max_1, bbox_req_stream_rsc_dat_x_min_1, bbox_req_stream_rsc_dat_z,
      bbox_req_stream_rsc_dat_y, bbox_req_stream_rsc_dat_x, bbox_req_stream_rsc_dat_d,
      bbox_req_stream_rsc_dat_d_1, bbox_req_stream_rsc_dat_d_2, bbox_req_stream_rsc_dat_d_3,
      bbox_req_stream_rsc_dat_d_4, bbox_req_stream_rsc_dat_d_5, bbox_req_stream_rsc_dat_d_6,
      bbox_req_stream_rsc_dat_d_7, bbox_req_stream_rsc_dat_rid, bbox_req_stream_rsc_vld,
      bbox_req_stream_rsc_rdy, ist_req_stream_rsc_dat_d, ist_req_stream_rsc_dat_d_1,
      ist_req_stream_rsc_dat_d_2, ist_req_stream_rsc_dat_d_3, ist_req_stream_rsc_dat_d_4,
      ist_req_stream_rsc_dat_d_5, ist_req_stream_rsc_dat_d_6, ist_req_stream_rsc_dat_d_7,
      ist_req_stream_rsc_dat_d_8, ist_req_stream_rsc_dat_d_9, ist_req_stream_rsc_dat_d_10,
      ist_req_stream_rsc_dat_d_11, ist_req_stream_rsc_dat_d_12, ist_req_stream_rsc_dat_d_13,
      ist_req_stream_rsc_dat_d_14, ist_req_stream_rsc_dat_d_15, ist_req_stream_rsc_dat_d_16,
      ist_req_stream_rsc_dat_rid, ist_req_stream_rsc_vld, ist_req_stream_rsc_rdy,
      trv_req_stream_rsc_dat_d, trv_req_stream_rsc_dat_d_1, trv_req_stream_rsc_dat_d_2,
      trv_req_stream_rsc_dat_d_3, trv_req_stream_rsc_dat_d_4, trv_req_stream_rsc_dat_d_5,
      trv_req_stream_rsc_dat_d_6, trv_req_stream_rsc_dat_d_7, trv_req_stream_rsc_dat_d_8,
      trv_req_stream_rsc_dat_d_9, trv_req_stream_rsc_dat_d_10, trv_req_stream_rsc_dat_d_11,
      trv_req_stream_rsc_dat_d_12, trv_req_stream_rsc_dat_d_13, trv_req_stream_rsc_dat_rid,
      trv_req_stream_rsc_vld, trv_req_stream_rsc_rdy, bbox_resp_stream_rsc_dat_left_first,
      bbox_resp_stream_rsc_dat_right_hit, bbox_resp_stream_rsc_dat_left_hit, bbox_resp_stream_rsc_dat_d,
      bbox_resp_stream_rsc_dat_d_1, bbox_resp_stream_rsc_dat_d_2, bbox_resp_stream_rsc_dat_d_3,
      bbox_resp_stream_rsc_dat_d_4, bbox_resp_stream_rsc_dat_d_5, bbox_resp_stream_rsc_dat_rid,
      bbox_resp_stream_rsc_vld, bbox_resp_stream_rsc_rdy, ist_resp_stream_rsc_dat_d,
      ist_resp_stream_rsc_dat_d_1, ist_resp_stream_rsc_dat_d_2, ist_resp_stream_rsc_dat_intersected,
      ist_resp_stream_rsc_dat_rid, ist_resp_stream_rsc_vld, ist_resp_stream_rsc_rdy
);
  input clk;
  input arst_n;
  input [31:0] init_req_stream_rsc_dat_d;
  input [31:0] init_req_stream_rsc_dat_d_1;
  input [31:0] init_req_stream_rsc_dat_d_2;
  input [31:0] init_req_stream_rsc_dat_d_3;
  input [31:0] init_req_stream_rsc_dat_d_4;
  input [31:0] init_req_stream_rsc_dat_d_5;
  input [31:0] init_req_stream_rsc_dat_d_6;
  input [31:0] init_req_stream_rsc_dat_d_7;
  input [31:0] init_req_stream_rsc_dat_d_8;
  input [31:0] init_req_stream_rsc_dat_d_9;
  input [31:0] init_req_stream_rsc_dat_d_10;
  input [9:0] init_req_stream_rsc_dat_rid;
  input init_req_stream_rsc_vld;
  output init_req_stream_rsc_rdy;
  input [7:0] bbox_req_stream_rsc_dat_z_max;
  input [7:0] bbox_req_stream_rsc_dat_z_min;
  input [7:0] bbox_req_stream_rsc_dat_y_max;
  input [7:0] bbox_req_stream_rsc_dat_y_min;
  input [7:0] bbox_req_stream_rsc_dat_x_max;
  input [7:0] bbox_req_stream_rsc_dat_x_min;
  input [7:0] bbox_req_stream_rsc_dat_z_max_1;
  input [7:0] bbox_req_stream_rsc_dat_z_min_1;
  input [7:0] bbox_req_stream_rsc_dat_y_max_1;
  input [7:0] bbox_req_stream_rsc_dat_y_min_1;
  input [7:0] bbox_req_stream_rsc_dat_x_max_1;
  input [7:0] bbox_req_stream_rsc_dat_x_min_1;
  input [7:0] bbox_req_stream_rsc_dat_z;
  input [7:0] bbox_req_stream_rsc_dat_y;
  input [7:0] bbox_req_stream_rsc_dat_x;
  input [31:0] bbox_req_stream_rsc_dat_d;
  input [31:0] bbox_req_stream_rsc_dat_d_1;
  input [31:0] bbox_req_stream_rsc_dat_d_2;
  input [31:0] bbox_req_stream_rsc_dat_d_3;
  input [31:0] bbox_req_stream_rsc_dat_d_4;
  input [31:0] bbox_req_stream_rsc_dat_d_5;
  input [31:0] bbox_req_stream_rsc_dat_d_6;
  input [31:0] bbox_req_stream_rsc_dat_d_7;
  input [9:0] bbox_req_stream_rsc_dat_rid;
  input bbox_req_stream_rsc_vld;
  output bbox_req_stream_rsc_rdy;
  input [31:0] ist_req_stream_rsc_dat_d;
  input [31:0] ist_req_stream_rsc_dat_d_1;
  input [31:0] ist_req_stream_rsc_dat_d_2;
  input [31:0] ist_req_stream_rsc_dat_d_3;
  input [31:0] ist_req_stream_rsc_dat_d_4;
  input [31:0] ist_req_stream_rsc_dat_d_5;
  input [31:0] ist_req_stream_rsc_dat_d_6;
  input [31:0] ist_req_stream_rsc_dat_d_7;
  input [31:0] ist_req_stream_rsc_dat_d_8;
  input [31:0] ist_req_stream_rsc_dat_d_9;
  input [31:0] ist_req_stream_rsc_dat_d_10;
  input [31:0] ist_req_stream_rsc_dat_d_11;
  input [31:0] ist_req_stream_rsc_dat_d_12;
  input [31:0] ist_req_stream_rsc_dat_d_13;
  input [31:0] ist_req_stream_rsc_dat_d_14;
  input [31:0] ist_req_stream_rsc_dat_d_15;
  input [31:0] ist_req_stream_rsc_dat_d_16;
  input [9:0] ist_req_stream_rsc_dat_rid;
  input ist_req_stream_rsc_vld;
  output ist_req_stream_rsc_rdy;
  output [31:0] trv_req_stream_rsc_dat_d;
  output [31:0] trv_req_stream_rsc_dat_d_1;
  output [31:0] trv_req_stream_rsc_dat_d_2;
  output [31:0] trv_req_stream_rsc_dat_d_3;
  output [31:0] trv_req_stream_rsc_dat_d_4;
  output [31:0] trv_req_stream_rsc_dat_d_5;
  output [31:0] trv_req_stream_rsc_dat_d_6;
  output [31:0] trv_req_stream_rsc_dat_d_7;
  output [31:0] trv_req_stream_rsc_dat_d_8;
  output [31:0] trv_req_stream_rsc_dat_d_9;
  output [31:0] trv_req_stream_rsc_dat_d_10;
  output [31:0] trv_req_stream_rsc_dat_d_11;
  output [31:0] trv_req_stream_rsc_dat_d_12;
  output [31:0] trv_req_stream_rsc_dat_d_13;
  output [9:0] trv_req_stream_rsc_dat_rid;
  output trv_req_stream_rsc_vld;
  input trv_req_stream_rsc_rdy;
  output bbox_resp_stream_rsc_dat_left_first;
  output bbox_resp_stream_rsc_dat_right_hit;
  output bbox_resp_stream_rsc_dat_left_hit;
  output [31:0] bbox_resp_stream_rsc_dat_d;
  output [31:0] bbox_resp_stream_rsc_dat_d_1;
  output [31:0] bbox_resp_stream_rsc_dat_d_2;
  output [31:0] bbox_resp_stream_rsc_dat_d_3;
  output [31:0] bbox_resp_stream_rsc_dat_d_4;
  output [31:0] bbox_resp_stream_rsc_dat_d_5;
  output [9:0] bbox_resp_stream_rsc_dat_rid;
  output bbox_resp_stream_rsc_vld;
  input bbox_resp_stream_rsc_rdy;
  output [31:0] ist_resp_stream_rsc_dat_d;
  output [31:0] ist_resp_stream_rsc_dat_d_1;
  output [31:0] ist_resp_stream_rsc_dat_d_2;
  output ist_resp_stream_rsc_dat_intersected;
  output [9:0] ist_resp_stream_rsc_dat_rid;
  output ist_resp_stream_rsc_vld;
  input ist_resp_stream_rsc_rdy;


  // Interconnect Declarations
  wire [457:0] trv_req_stream_rsc_dat_n_init_inst;
  wire [204:0] bbox_resp_stream_rsc_dat_n_bbox_inst;
  wire [106:0] ist_resp_stream_rsc_dat_n_ist_inst;
  wire init_req_stream_rsc_rdy_n_init_inst_bud;
  wire trv_req_stream_rsc_vld_n_init_inst_bud;
  wire bbox_req_stream_rsc_rdy_n_bbox_inst_bud;
  wire bbox_resp_stream_rsc_vld_n_bbox_inst_bud;
  wire ist_req_stream_rsc_rdy_n_ist_inst_bud;
  wire ist_resp_stream_rsc_vld_n_ist_inst_bud;


  // Interconnect Declarations for Component Instantiations 
  wire [361:0] nl_init_inst_init_req_stream_rsc_dat;
  assign nl_init_inst_init_req_stream_rsc_dat = {init_req_stream_rsc_dat_d , init_req_stream_rsc_dat_d_1
      , init_req_stream_rsc_dat_d_2 , init_req_stream_rsc_dat_d_3 , init_req_stream_rsc_dat_d_4
      , init_req_stream_rsc_dat_d_5 , init_req_stream_rsc_dat_d_6 , init_req_stream_rsc_dat_d_7
      , init_req_stream_rsc_dat_d_8 , init_req_stream_rsc_dat_d_9 , init_req_stream_rsc_dat_d_10
      , init_req_stream_rsc_dat_rid};
  wire [385:0] nl_bbox_inst_bbox_req_stream_rsc_dat;
  assign nl_bbox_inst_bbox_req_stream_rsc_dat = {bbox_req_stream_rsc_dat_z_max ,
      bbox_req_stream_rsc_dat_z_min , bbox_req_stream_rsc_dat_y_max , bbox_req_stream_rsc_dat_y_min
      , bbox_req_stream_rsc_dat_x_max , bbox_req_stream_rsc_dat_x_min , bbox_req_stream_rsc_dat_z_max_1
      , bbox_req_stream_rsc_dat_z_min_1 , bbox_req_stream_rsc_dat_y_max_1 , bbox_req_stream_rsc_dat_y_min_1
      , bbox_req_stream_rsc_dat_x_max_1 , bbox_req_stream_rsc_dat_x_min_1 , bbox_req_stream_rsc_dat_z
      , bbox_req_stream_rsc_dat_y , bbox_req_stream_rsc_dat_x , bbox_req_stream_rsc_dat_d
      , bbox_req_stream_rsc_dat_d_1 , bbox_req_stream_rsc_dat_d_2 , bbox_req_stream_rsc_dat_d_3
      , bbox_req_stream_rsc_dat_d_4 , bbox_req_stream_rsc_dat_d_5 , bbox_req_stream_rsc_dat_d_6
      , bbox_req_stream_rsc_dat_d_7 , bbox_req_stream_rsc_dat_rid};
  wire [553:0] nl_ist_inst_ist_req_stream_rsc_dat;
  assign nl_ist_inst_ist_req_stream_rsc_dat = {ist_req_stream_rsc_dat_d , ist_req_stream_rsc_dat_d_1
      , ist_req_stream_rsc_dat_d_2 , ist_req_stream_rsc_dat_d_3 , ist_req_stream_rsc_dat_d_4
      , ist_req_stream_rsc_dat_d_5 , ist_req_stream_rsc_dat_d_6 , ist_req_stream_rsc_dat_d_7
      , ist_req_stream_rsc_dat_d_8 , ist_req_stream_rsc_dat_d_9 , ist_req_stream_rsc_dat_d_10
      , ist_req_stream_rsc_dat_d_11 , ist_req_stream_rsc_dat_d_12 , ist_req_stream_rsc_dat_d_13
      , ist_req_stream_rsc_dat_d_14 , ist_req_stream_rsc_dat_d_15 , ist_req_stream_rsc_dat_d_16
      , ist_req_stream_rsc_dat_rid};
  init init_inst (
      .clk(clk),
      .arst_n(arst_n),
      .init_req_stream_rsc_dat(nl_init_inst_init_req_stream_rsc_dat[361:0]),
      .init_req_stream_rsc_vld(init_req_stream_rsc_vld),
      .init_req_stream_rsc_rdy(init_req_stream_rsc_rdy_n_init_inst_bud),
      .trv_req_stream_rsc_dat(trv_req_stream_rsc_dat_n_init_inst),
      .trv_req_stream_rsc_vld(trv_req_stream_rsc_vld_n_init_inst_bud),
      .trv_req_stream_rsc_rdy(trv_req_stream_rsc_rdy)
    );
  bbox bbox_inst (
      .clk(clk),
      .arst_n(arst_n),
      .bbox_req_stream_rsc_dat(nl_bbox_inst_bbox_req_stream_rsc_dat[385:0]),
      .bbox_req_stream_rsc_vld(bbox_req_stream_rsc_vld),
      .bbox_req_stream_rsc_rdy(bbox_req_stream_rsc_rdy_n_bbox_inst_bud),
      .bbox_resp_stream_rsc_dat(bbox_resp_stream_rsc_dat_n_bbox_inst),
      .bbox_resp_stream_rsc_vld(bbox_resp_stream_rsc_vld_n_bbox_inst_bud),
      .bbox_resp_stream_rsc_rdy(bbox_resp_stream_rsc_rdy)
    );
  ist ist_inst (
      .clk(clk),
      .arst_n(arst_n),
      .ist_req_stream_rsc_dat(nl_ist_inst_ist_req_stream_rsc_dat[553:0]),
      .ist_req_stream_rsc_vld(ist_req_stream_rsc_vld),
      .ist_req_stream_rsc_rdy(ist_req_stream_rsc_rdy_n_ist_inst_bud),
      .ist_resp_stream_rsc_dat(ist_resp_stream_rsc_dat_n_ist_inst),
      .ist_resp_stream_rsc_vld(ist_resp_stream_rsc_vld_n_ist_inst_bud),
      .ist_resp_stream_rsc_rdy(ist_resp_stream_rsc_rdy)
    );
  assign init_req_stream_rsc_rdy = init_req_stream_rsc_rdy_n_init_inst_bud;
  assign trv_req_stream_rsc_dat_rid = trv_req_stream_rsc_dat_n_init_inst[9:0];
  assign trv_req_stream_rsc_dat_d_13 = trv_req_stream_rsc_dat_n_init_inst[41:10];
  assign trv_req_stream_rsc_dat_d_12 = trv_req_stream_rsc_dat_n_init_inst[73:42];
  assign trv_req_stream_rsc_dat_d_11 = trv_req_stream_rsc_dat_n_init_inst[105:74];
  assign trv_req_stream_rsc_dat_d_10 = trv_req_stream_rsc_dat_n_init_inst[137:106];
  assign trv_req_stream_rsc_dat_d_9 = trv_req_stream_rsc_dat_n_init_inst[169:138];
  assign trv_req_stream_rsc_dat_d_8 = trv_req_stream_rsc_dat_n_init_inst[201:170];
  assign trv_req_stream_rsc_dat_d_7 = trv_req_stream_rsc_dat_n_init_inst[233:202];
  assign trv_req_stream_rsc_dat_d_6 = trv_req_stream_rsc_dat_n_init_inst[265:234];
  assign trv_req_stream_rsc_dat_d_5 = trv_req_stream_rsc_dat_n_init_inst[297:266];
  assign trv_req_stream_rsc_dat_d_4 = trv_req_stream_rsc_dat_n_init_inst[329:298];
  assign trv_req_stream_rsc_dat_d_3 = trv_req_stream_rsc_dat_n_init_inst[361:330];
  assign trv_req_stream_rsc_dat_d_2 = trv_req_stream_rsc_dat_n_init_inst[393:362];
  assign trv_req_stream_rsc_dat_d_1 = trv_req_stream_rsc_dat_n_init_inst[425:394];
  assign trv_req_stream_rsc_dat_d = trv_req_stream_rsc_dat_n_init_inst[457:426];
  assign bbox_resp_stream_rsc_dat_rid = bbox_resp_stream_rsc_dat_n_bbox_inst[9:0];
  assign bbox_resp_stream_rsc_dat_d_5 = bbox_resp_stream_rsc_dat_n_bbox_inst[41:10];
  assign bbox_resp_stream_rsc_dat_d_4 = bbox_resp_stream_rsc_dat_n_bbox_inst[73:42];
  assign bbox_resp_stream_rsc_dat_d_3 = bbox_resp_stream_rsc_dat_n_bbox_inst[105:74];
  assign bbox_resp_stream_rsc_dat_d_2 = bbox_resp_stream_rsc_dat_n_bbox_inst[137:106];
  assign bbox_resp_stream_rsc_dat_d_1 = bbox_resp_stream_rsc_dat_n_bbox_inst[169:138];
  assign bbox_resp_stream_rsc_dat_d = bbox_resp_stream_rsc_dat_n_bbox_inst[201:170];
  assign bbox_resp_stream_rsc_dat_left_hit = bbox_resp_stream_rsc_dat_n_bbox_inst[202];
  assign bbox_resp_stream_rsc_dat_right_hit = bbox_resp_stream_rsc_dat_n_bbox_inst[203];
  assign bbox_resp_stream_rsc_dat_left_first = bbox_resp_stream_rsc_dat_n_bbox_inst[204];
  assign ist_resp_stream_rsc_dat_rid = ist_resp_stream_rsc_dat_n_ist_inst[9:0];
  assign ist_resp_stream_rsc_dat_intersected = ist_resp_stream_rsc_dat_n_ist_inst[10];
  assign ist_resp_stream_rsc_dat_d_2 = ist_resp_stream_rsc_dat_n_ist_inst[42:11];
  assign ist_resp_stream_rsc_dat_d_1 = ist_resp_stream_rsc_dat_n_ist_inst[74:43];
  assign ist_resp_stream_rsc_dat_d = ist_resp_stream_rsc_dat_n_ist_inst[106:75];
  assign bbox_req_stream_rsc_rdy = bbox_req_stream_rsc_rdy_n_bbox_inst_bud;
  assign ist_req_stream_rsc_rdy = ist_req_stream_rsc_rdy_n_ist_inst_bud;
  assign trv_req_stream_rsc_vld = trv_req_stream_rsc_vld_n_init_inst_bud;
  assign bbox_resp_stream_rsc_vld = bbox_resp_stream_rsc_vld_n_bbox_inst_bud;
  assign ist_resp_stream_rsc_vld = ist_resp_stream_rsc_vld_n_ist_inst_bud;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    rtcore
// ------------------------------------------------------------------


module rtcore (
  clk, arst_n, init_req_stream_rsc_dat, init_req_stream_rsc_vld, init_req_stream_rsc_rdy,
      bbox_req_stream_rsc_dat, bbox_req_stream_rsc_vld, bbox_req_stream_rsc_rdy,
      ist_req_stream_rsc_dat, ist_req_stream_rsc_vld, ist_req_stream_rsc_rdy, trv_req_stream_rsc_dat,
      trv_req_stream_rsc_vld, trv_req_stream_rsc_rdy, bbox_resp_stream_rsc_dat, bbox_resp_stream_rsc_vld,
      bbox_resp_stream_rsc_rdy, ist_resp_stream_rsc_dat, ist_resp_stream_rsc_vld,
      ist_resp_stream_rsc_rdy
);
  input clk;
  input arst_n;
  input [361:0] init_req_stream_rsc_dat;
  input init_req_stream_rsc_vld;
  output init_req_stream_rsc_rdy;
  input [385:0] bbox_req_stream_rsc_dat;
  input bbox_req_stream_rsc_vld;
  output bbox_req_stream_rsc_rdy;
  input [553:0] ist_req_stream_rsc_dat;
  input ist_req_stream_rsc_vld;
  output ist_req_stream_rsc_rdy;
  output [457:0] trv_req_stream_rsc_dat;
  output trv_req_stream_rsc_vld;
  input trv_req_stream_rsc_rdy;
  output [204:0] bbox_resp_stream_rsc_dat;
  output bbox_resp_stream_rsc_vld;
  input bbox_resp_stream_rsc_rdy;
  output [106:0] ist_resp_stream_rsc_dat;
  output ist_resp_stream_rsc_vld;
  input ist_resp_stream_rsc_rdy;


  // Interconnect Declarations
  wire [31:0] trv_req_stream_rsc_dat_d;
  wire [31:0] trv_req_stream_rsc_dat_d_1;
  wire [31:0] trv_req_stream_rsc_dat_d_2;
  wire [31:0] trv_req_stream_rsc_dat_d_3;
  wire [31:0] trv_req_stream_rsc_dat_d_4;
  wire [31:0] trv_req_stream_rsc_dat_d_5;
  wire [31:0] trv_req_stream_rsc_dat_d_6;
  wire [31:0] trv_req_stream_rsc_dat_d_7;
  wire [31:0] trv_req_stream_rsc_dat_d_8;
  wire [31:0] trv_req_stream_rsc_dat_d_9;
  wire [31:0] trv_req_stream_rsc_dat_d_10;
  wire [31:0] trv_req_stream_rsc_dat_d_11;
  wire [31:0] trv_req_stream_rsc_dat_d_12;
  wire [31:0] trv_req_stream_rsc_dat_d_13;
  wire [9:0] trv_req_stream_rsc_dat_rid;
  wire bbox_resp_stream_rsc_dat_left_first;
  wire bbox_resp_stream_rsc_dat_right_hit;
  wire bbox_resp_stream_rsc_dat_left_hit;
  wire [31:0] bbox_resp_stream_rsc_dat_d;
  wire [31:0] bbox_resp_stream_rsc_dat_d_1;
  wire [31:0] bbox_resp_stream_rsc_dat_d_2;
  wire [31:0] bbox_resp_stream_rsc_dat_d_3;
  wire [31:0] bbox_resp_stream_rsc_dat_d_4;
  wire [31:0] bbox_resp_stream_rsc_dat_d_5;
  wire [9:0] bbox_resp_stream_rsc_dat_rid;
  wire [31:0] ist_resp_stream_rsc_dat_d;
  wire [31:0] ist_resp_stream_rsc_dat_d_1;
  wire [31:0] ist_resp_stream_rsc_dat_d_2;
  wire ist_resp_stream_rsc_dat_intersected;
  wire [9:0] ist_resp_stream_rsc_dat_rid;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_rtcore_struct_inst_init_req_stream_rsc_dat_d;
  assign nl_rtcore_struct_inst_init_req_stream_rsc_dat_d = init_req_stream_rsc_dat[361:330];
  wire [31:0] nl_rtcore_struct_inst_init_req_stream_rsc_dat_d_1;
  assign nl_rtcore_struct_inst_init_req_stream_rsc_dat_d_1 = init_req_stream_rsc_dat[329:298];
  wire [31:0] nl_rtcore_struct_inst_init_req_stream_rsc_dat_d_2;
  assign nl_rtcore_struct_inst_init_req_stream_rsc_dat_d_2 = init_req_stream_rsc_dat[297:266];
  wire [31:0] nl_rtcore_struct_inst_init_req_stream_rsc_dat_d_3;
  assign nl_rtcore_struct_inst_init_req_stream_rsc_dat_d_3 = init_req_stream_rsc_dat[265:234];
  wire [31:0] nl_rtcore_struct_inst_init_req_stream_rsc_dat_d_4;
  assign nl_rtcore_struct_inst_init_req_stream_rsc_dat_d_4 = init_req_stream_rsc_dat[233:202];
  wire [31:0] nl_rtcore_struct_inst_init_req_stream_rsc_dat_d_5;
  assign nl_rtcore_struct_inst_init_req_stream_rsc_dat_d_5 = init_req_stream_rsc_dat[201:170];
  wire [31:0] nl_rtcore_struct_inst_init_req_stream_rsc_dat_d_6;
  assign nl_rtcore_struct_inst_init_req_stream_rsc_dat_d_6 = init_req_stream_rsc_dat[169:138];
  wire [31:0] nl_rtcore_struct_inst_init_req_stream_rsc_dat_d_7;
  assign nl_rtcore_struct_inst_init_req_stream_rsc_dat_d_7 = init_req_stream_rsc_dat[137:106];
  wire [31:0] nl_rtcore_struct_inst_init_req_stream_rsc_dat_d_8;
  assign nl_rtcore_struct_inst_init_req_stream_rsc_dat_d_8 = init_req_stream_rsc_dat[105:74];
  wire [31:0] nl_rtcore_struct_inst_init_req_stream_rsc_dat_d_9;
  assign nl_rtcore_struct_inst_init_req_stream_rsc_dat_d_9 = init_req_stream_rsc_dat[73:42];
  wire [31:0] nl_rtcore_struct_inst_init_req_stream_rsc_dat_d_10;
  assign nl_rtcore_struct_inst_init_req_stream_rsc_dat_d_10 = init_req_stream_rsc_dat[41:10];
  wire [9:0] nl_rtcore_struct_inst_init_req_stream_rsc_dat_rid;
  assign nl_rtcore_struct_inst_init_req_stream_rsc_dat_rid = init_req_stream_rsc_dat[9:0];
  wire [7:0] nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_z_max;
  assign nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_z_max = bbox_req_stream_rsc_dat[385:378];
  wire [7:0] nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_z_min;
  assign nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_z_min = bbox_req_stream_rsc_dat[377:370];
  wire [7:0] nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_y_max;
  assign nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_y_max = bbox_req_stream_rsc_dat[369:362];
  wire [7:0] nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_y_min;
  assign nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_y_min = bbox_req_stream_rsc_dat[361:354];
  wire [7:0] nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_x_max;
  assign nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_x_max = bbox_req_stream_rsc_dat[353:346];
  wire [7:0] nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_x_min;
  assign nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_x_min = bbox_req_stream_rsc_dat[345:338];
  wire [7:0] nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_z_max_1;
  assign nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_z_max_1 = bbox_req_stream_rsc_dat[337:330];
  wire [7:0] nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_z_min_1;
  assign nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_z_min_1 = bbox_req_stream_rsc_dat[329:322];
  wire [7:0] nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_y_max_1;
  assign nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_y_max_1 = bbox_req_stream_rsc_dat[321:314];
  wire [7:0] nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_y_min_1;
  assign nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_y_min_1 = bbox_req_stream_rsc_dat[313:306];
  wire [7:0] nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_x_max_1;
  assign nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_x_max_1 = bbox_req_stream_rsc_dat[305:298];
  wire [7:0] nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_x_min_1;
  assign nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_x_min_1 = bbox_req_stream_rsc_dat[297:290];
  wire [7:0] nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_z;
  assign nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_z = bbox_req_stream_rsc_dat[289:282];
  wire [7:0] nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_y;
  assign nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_y = bbox_req_stream_rsc_dat[281:274];
  wire [7:0] nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_x;
  assign nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_x = bbox_req_stream_rsc_dat[273:266];
  wire [31:0] nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_d;
  assign nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_d = bbox_req_stream_rsc_dat[265:234];
  wire [31:0] nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_d_1;
  assign nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_d_1 = bbox_req_stream_rsc_dat[233:202];
  wire [31:0] nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_d_2;
  assign nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_d_2 = bbox_req_stream_rsc_dat[201:170];
  wire [31:0] nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_d_3;
  assign nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_d_3 = bbox_req_stream_rsc_dat[169:138];
  wire [31:0] nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_d_4;
  assign nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_d_4 = bbox_req_stream_rsc_dat[137:106];
  wire [31:0] nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_d_5;
  assign nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_d_5 = bbox_req_stream_rsc_dat[105:74];
  wire [31:0] nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_d_6;
  assign nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_d_6 = bbox_req_stream_rsc_dat[73:42];
  wire [31:0] nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_d_7;
  assign nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_d_7 = bbox_req_stream_rsc_dat[41:10];
  wire [9:0] nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_rid;
  assign nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_rid = bbox_req_stream_rsc_dat[9:0];
  wire [31:0] nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d;
  assign nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d = ist_req_stream_rsc_dat[553:522];
  wire [31:0] nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_1;
  assign nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_1 = ist_req_stream_rsc_dat[521:490];
  wire [31:0] nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_2;
  assign nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_2 = ist_req_stream_rsc_dat[489:458];
  wire [31:0] nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_3;
  assign nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_3 = ist_req_stream_rsc_dat[457:426];
  wire [31:0] nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_4;
  assign nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_4 = ist_req_stream_rsc_dat[425:394];
  wire [31:0] nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_5;
  assign nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_5 = ist_req_stream_rsc_dat[393:362];
  wire [31:0] nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_6;
  assign nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_6 = ist_req_stream_rsc_dat[361:330];
  wire [31:0] nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_7;
  assign nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_7 = ist_req_stream_rsc_dat[329:298];
  wire [31:0] nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_8;
  assign nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_8 = ist_req_stream_rsc_dat[297:266];
  wire [31:0] nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_9;
  assign nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_9 = ist_req_stream_rsc_dat[265:234];
  wire [31:0] nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_10;
  assign nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_10 = ist_req_stream_rsc_dat[233:202];
  wire [31:0] nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_11;
  assign nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_11 = ist_req_stream_rsc_dat[201:170];
  wire [31:0] nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_12;
  assign nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_12 = ist_req_stream_rsc_dat[169:138];
  wire [31:0] nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_13;
  assign nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_13 = ist_req_stream_rsc_dat[137:106];
  wire [31:0] nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_14;
  assign nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_14 = ist_req_stream_rsc_dat[105:74];
  wire [31:0] nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_15;
  assign nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_15 = ist_req_stream_rsc_dat[73:42];
  wire [31:0] nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_16;
  assign nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_16 = ist_req_stream_rsc_dat[41:10];
  wire [9:0] nl_rtcore_struct_inst_ist_req_stream_rsc_dat_rid;
  assign nl_rtcore_struct_inst_ist_req_stream_rsc_dat_rid = ist_req_stream_rsc_dat[9:0];
  rtcore_struct rtcore_struct_inst (
      .clk(clk),
      .arst_n(arst_n),
      .init_req_stream_rsc_dat_d(nl_rtcore_struct_inst_init_req_stream_rsc_dat_d[31:0]),
      .init_req_stream_rsc_dat_d_1(nl_rtcore_struct_inst_init_req_stream_rsc_dat_d_1[31:0]),
      .init_req_stream_rsc_dat_d_2(nl_rtcore_struct_inst_init_req_stream_rsc_dat_d_2[31:0]),
      .init_req_stream_rsc_dat_d_3(nl_rtcore_struct_inst_init_req_stream_rsc_dat_d_3[31:0]),
      .init_req_stream_rsc_dat_d_4(nl_rtcore_struct_inst_init_req_stream_rsc_dat_d_4[31:0]),
      .init_req_stream_rsc_dat_d_5(nl_rtcore_struct_inst_init_req_stream_rsc_dat_d_5[31:0]),
      .init_req_stream_rsc_dat_d_6(nl_rtcore_struct_inst_init_req_stream_rsc_dat_d_6[31:0]),
      .init_req_stream_rsc_dat_d_7(nl_rtcore_struct_inst_init_req_stream_rsc_dat_d_7[31:0]),
      .init_req_stream_rsc_dat_d_8(nl_rtcore_struct_inst_init_req_stream_rsc_dat_d_8[31:0]),
      .init_req_stream_rsc_dat_d_9(nl_rtcore_struct_inst_init_req_stream_rsc_dat_d_9[31:0]),
      .init_req_stream_rsc_dat_d_10(nl_rtcore_struct_inst_init_req_stream_rsc_dat_d_10[31:0]),
      .init_req_stream_rsc_dat_rid(nl_rtcore_struct_inst_init_req_stream_rsc_dat_rid[9:0]),
      .init_req_stream_rsc_vld(init_req_stream_rsc_vld),
      .init_req_stream_rsc_rdy(init_req_stream_rsc_rdy),
      .bbox_req_stream_rsc_dat_z_max(nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_z_max[7:0]),
      .bbox_req_stream_rsc_dat_z_min(nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_z_min[7:0]),
      .bbox_req_stream_rsc_dat_y_max(nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_y_max[7:0]),
      .bbox_req_stream_rsc_dat_y_min(nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_y_min[7:0]),
      .bbox_req_stream_rsc_dat_x_max(nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_x_max[7:0]),
      .bbox_req_stream_rsc_dat_x_min(nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_x_min[7:0]),
      .bbox_req_stream_rsc_dat_z_max_1(nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_z_max_1[7:0]),
      .bbox_req_stream_rsc_dat_z_min_1(nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_z_min_1[7:0]),
      .bbox_req_stream_rsc_dat_y_max_1(nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_y_max_1[7:0]),
      .bbox_req_stream_rsc_dat_y_min_1(nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_y_min_1[7:0]),
      .bbox_req_stream_rsc_dat_x_max_1(nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_x_max_1[7:0]),
      .bbox_req_stream_rsc_dat_x_min_1(nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_x_min_1[7:0]),
      .bbox_req_stream_rsc_dat_z(nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_z[7:0]),
      .bbox_req_stream_rsc_dat_y(nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_y[7:0]),
      .bbox_req_stream_rsc_dat_x(nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_x[7:0]),
      .bbox_req_stream_rsc_dat_d(nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_d[31:0]),
      .bbox_req_stream_rsc_dat_d_1(nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_d_1[31:0]),
      .bbox_req_stream_rsc_dat_d_2(nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_d_2[31:0]),
      .bbox_req_stream_rsc_dat_d_3(nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_d_3[31:0]),
      .bbox_req_stream_rsc_dat_d_4(nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_d_4[31:0]),
      .bbox_req_stream_rsc_dat_d_5(nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_d_5[31:0]),
      .bbox_req_stream_rsc_dat_d_6(nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_d_6[31:0]),
      .bbox_req_stream_rsc_dat_d_7(nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_d_7[31:0]),
      .bbox_req_stream_rsc_dat_rid(nl_rtcore_struct_inst_bbox_req_stream_rsc_dat_rid[9:0]),
      .bbox_req_stream_rsc_vld(bbox_req_stream_rsc_vld),
      .bbox_req_stream_rsc_rdy(bbox_req_stream_rsc_rdy),
      .ist_req_stream_rsc_dat_d(nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d[31:0]),
      .ist_req_stream_rsc_dat_d_1(nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_1[31:0]),
      .ist_req_stream_rsc_dat_d_2(nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_2[31:0]),
      .ist_req_stream_rsc_dat_d_3(nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_3[31:0]),
      .ist_req_stream_rsc_dat_d_4(nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_4[31:0]),
      .ist_req_stream_rsc_dat_d_5(nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_5[31:0]),
      .ist_req_stream_rsc_dat_d_6(nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_6[31:0]),
      .ist_req_stream_rsc_dat_d_7(nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_7[31:0]),
      .ist_req_stream_rsc_dat_d_8(nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_8[31:0]),
      .ist_req_stream_rsc_dat_d_9(nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_9[31:0]),
      .ist_req_stream_rsc_dat_d_10(nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_10[31:0]),
      .ist_req_stream_rsc_dat_d_11(nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_11[31:0]),
      .ist_req_stream_rsc_dat_d_12(nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_12[31:0]),
      .ist_req_stream_rsc_dat_d_13(nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_13[31:0]),
      .ist_req_stream_rsc_dat_d_14(nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_14[31:0]),
      .ist_req_stream_rsc_dat_d_15(nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_15[31:0]),
      .ist_req_stream_rsc_dat_d_16(nl_rtcore_struct_inst_ist_req_stream_rsc_dat_d_16[31:0]),
      .ist_req_stream_rsc_dat_rid(nl_rtcore_struct_inst_ist_req_stream_rsc_dat_rid[9:0]),
      .ist_req_stream_rsc_vld(ist_req_stream_rsc_vld),
      .ist_req_stream_rsc_rdy(ist_req_stream_rsc_rdy),
      .trv_req_stream_rsc_dat_d(trv_req_stream_rsc_dat_d),
      .trv_req_stream_rsc_dat_d_1(trv_req_stream_rsc_dat_d_1),
      .trv_req_stream_rsc_dat_d_2(trv_req_stream_rsc_dat_d_2),
      .trv_req_stream_rsc_dat_d_3(trv_req_stream_rsc_dat_d_3),
      .trv_req_stream_rsc_dat_d_4(trv_req_stream_rsc_dat_d_4),
      .trv_req_stream_rsc_dat_d_5(trv_req_stream_rsc_dat_d_5),
      .trv_req_stream_rsc_dat_d_6(trv_req_stream_rsc_dat_d_6),
      .trv_req_stream_rsc_dat_d_7(trv_req_stream_rsc_dat_d_7),
      .trv_req_stream_rsc_dat_d_8(trv_req_stream_rsc_dat_d_8),
      .trv_req_stream_rsc_dat_d_9(trv_req_stream_rsc_dat_d_9),
      .trv_req_stream_rsc_dat_d_10(trv_req_stream_rsc_dat_d_10),
      .trv_req_stream_rsc_dat_d_11(trv_req_stream_rsc_dat_d_11),
      .trv_req_stream_rsc_dat_d_12(trv_req_stream_rsc_dat_d_12),
      .trv_req_stream_rsc_dat_d_13(trv_req_stream_rsc_dat_d_13),
      .trv_req_stream_rsc_dat_rid(trv_req_stream_rsc_dat_rid),
      .trv_req_stream_rsc_vld(trv_req_stream_rsc_vld),
      .trv_req_stream_rsc_rdy(trv_req_stream_rsc_rdy),
      .bbox_resp_stream_rsc_dat_left_first(bbox_resp_stream_rsc_dat_left_first),
      .bbox_resp_stream_rsc_dat_right_hit(bbox_resp_stream_rsc_dat_right_hit),
      .bbox_resp_stream_rsc_dat_left_hit(bbox_resp_stream_rsc_dat_left_hit),
      .bbox_resp_stream_rsc_dat_d(bbox_resp_stream_rsc_dat_d),
      .bbox_resp_stream_rsc_dat_d_1(bbox_resp_stream_rsc_dat_d_1),
      .bbox_resp_stream_rsc_dat_d_2(bbox_resp_stream_rsc_dat_d_2),
      .bbox_resp_stream_rsc_dat_d_3(bbox_resp_stream_rsc_dat_d_3),
      .bbox_resp_stream_rsc_dat_d_4(bbox_resp_stream_rsc_dat_d_4),
      .bbox_resp_stream_rsc_dat_d_5(bbox_resp_stream_rsc_dat_d_5),
      .bbox_resp_stream_rsc_dat_rid(bbox_resp_stream_rsc_dat_rid),
      .bbox_resp_stream_rsc_vld(bbox_resp_stream_rsc_vld),
      .bbox_resp_stream_rsc_rdy(bbox_resp_stream_rsc_rdy),
      .ist_resp_stream_rsc_dat_d(ist_resp_stream_rsc_dat_d),
      .ist_resp_stream_rsc_dat_d_1(ist_resp_stream_rsc_dat_d_1),
      .ist_resp_stream_rsc_dat_d_2(ist_resp_stream_rsc_dat_d_2),
      .ist_resp_stream_rsc_dat_intersected(ist_resp_stream_rsc_dat_intersected),
      .ist_resp_stream_rsc_dat_rid(ist_resp_stream_rsc_dat_rid),
      .ist_resp_stream_rsc_vld(ist_resp_stream_rsc_vld),
      .ist_resp_stream_rsc_rdy(ist_resp_stream_rsc_rdy)
    );
  assign trv_req_stream_rsc_dat = {trv_req_stream_rsc_dat_d , trv_req_stream_rsc_dat_d_1
      , trv_req_stream_rsc_dat_d_2 , trv_req_stream_rsc_dat_d_3 , trv_req_stream_rsc_dat_d_4
      , trv_req_stream_rsc_dat_d_5 , trv_req_stream_rsc_dat_d_6 , trv_req_stream_rsc_dat_d_7
      , trv_req_stream_rsc_dat_d_8 , trv_req_stream_rsc_dat_d_9 , trv_req_stream_rsc_dat_d_10
      , trv_req_stream_rsc_dat_d_11 , trv_req_stream_rsc_dat_d_12 , trv_req_stream_rsc_dat_d_13
      , trv_req_stream_rsc_dat_rid};
  assign bbox_resp_stream_rsc_dat = {bbox_resp_stream_rsc_dat_left_first , bbox_resp_stream_rsc_dat_right_hit
      , bbox_resp_stream_rsc_dat_left_hit , bbox_resp_stream_rsc_dat_d , bbox_resp_stream_rsc_dat_d_1
      , bbox_resp_stream_rsc_dat_d_2 , bbox_resp_stream_rsc_dat_d_3 , bbox_resp_stream_rsc_dat_d_4
      , bbox_resp_stream_rsc_dat_d_5 , bbox_resp_stream_rsc_dat_rid};
  assign ist_resp_stream_rsc_dat = {ist_resp_stream_rsc_dat_d , ist_resp_stream_rsc_dat_d_1
      , ist_resp_stream_rsc_dat_d_2 , ist_resp_stream_rsc_dat_intersected , ist_resp_stream_rsc_dat_rid};
endmodule



